magic
tech scmos
timestamp
<< pdiffusion >>
rect 420 440 421 441
rect 422 440 423 441
rect 423 440 424 441
rect 425 440 426 441
rect 420 441 426 445
rect 420 445 421 446
rect 422 445 423 446
rect 423 445 424 446
rect 425 445 426 446
rect 360 280 361 281
rect 362 280 363 281
rect 363 280 364 281
rect 365 280 366 281
rect 360 281 366 285
rect 360 285 361 286
rect 362 285 363 286
rect 363 285 364 286
rect 365 285 366 286
rect 80 480 81 481
rect 82 480 83 481
rect 83 480 84 481
rect 85 480 86 481
rect 80 481 86 485
rect 80 485 81 486
rect 82 485 83 486
rect 83 485 84 486
rect 85 485 86 486
rect 120 160 121 161
rect 122 160 123 161
rect 123 160 124 161
rect 125 160 126 161
rect 120 161 126 165
rect 120 165 121 166
rect 122 165 123 166
rect 123 165 124 166
rect 125 165 126 166
rect 460 580 461 581
rect 462 580 463 581
rect 463 580 464 581
rect 465 580 466 581
rect 460 581 466 585
rect 460 585 461 586
rect 462 585 463 586
rect 463 585 464 586
rect 465 585 466 586
rect 420 160 421 161
rect 422 160 423 161
rect 423 160 424 161
rect 425 160 426 161
rect 420 161 426 165
rect 420 165 421 166
rect 422 165 423 166
rect 423 165 424 166
rect 425 165 426 166
rect 520 20 521 21
rect 522 20 523 21
rect 523 20 524 21
rect 525 20 526 21
rect 520 21 526 25
rect 520 25 521 26
rect 522 25 523 26
rect 523 25 524 26
rect 525 25 526 26
rect 480 440 481 441
rect 482 440 483 441
rect 483 440 484 441
rect 485 440 486 441
rect 480 441 486 445
rect 480 445 481 446
rect 482 445 483 446
rect 483 445 484 446
rect 485 445 486 446
rect 500 180 501 181
rect 502 180 503 181
rect 503 180 504 181
rect 505 180 506 181
rect 500 181 506 185
rect 500 185 501 186
rect 502 185 503 186
rect 503 185 504 186
rect 505 185 506 186
rect 380 100 381 101
rect 382 100 383 101
rect 383 100 384 101
rect 385 100 386 101
rect 380 101 386 105
rect 380 105 381 106
rect 382 105 383 106
rect 383 105 384 106
rect 385 105 386 106
rect 580 280 581 281
rect 582 280 583 281
rect 583 280 584 281
rect 585 280 586 281
rect 580 281 586 285
rect 580 285 581 286
rect 582 285 583 286
rect 583 285 584 286
rect 585 285 586 286
rect 600 240 601 241
rect 602 240 603 241
rect 603 240 604 241
rect 605 240 606 241
rect 600 241 606 245
rect 600 245 601 246
rect 602 245 603 246
rect 603 245 604 246
rect 605 245 606 246
rect 320 160 321 161
rect 322 160 323 161
rect 323 160 324 161
rect 325 160 326 161
rect 320 161 326 165
rect 320 165 321 166
rect 322 165 323 166
rect 323 165 324 166
rect 325 165 326 166
rect 340 460 341 461
rect 342 460 343 461
rect 343 460 344 461
rect 345 460 346 461
rect 340 461 346 465
rect 340 465 341 466
rect 342 465 343 466
rect 343 465 344 466
rect 345 465 346 466
rect 40 280 41 281
rect 42 280 43 281
rect 43 280 44 281
rect 45 280 46 281
rect 40 281 46 285
rect 40 285 41 286
rect 42 285 43 286
rect 43 285 44 286
rect 45 285 46 286
rect 260 500 261 501
rect 262 500 263 501
rect 263 500 264 501
rect 265 500 266 501
rect 260 501 266 505
rect 260 505 261 506
rect 262 505 263 506
rect 263 505 264 506
rect 265 505 266 506
rect 480 360 481 361
rect 482 360 483 361
rect 483 360 484 361
rect 485 360 486 361
rect 480 361 486 365
rect 480 365 481 366
rect 482 365 483 366
rect 483 365 484 366
rect 485 365 486 366
rect 440 320 441 321
rect 442 320 443 321
rect 443 320 444 321
rect 445 320 446 321
rect 440 321 446 325
rect 440 325 441 326
rect 442 325 443 326
rect 443 325 444 326
rect 445 325 446 326
rect 280 60 281 61
rect 282 60 283 61
rect 283 60 284 61
rect 285 60 286 61
rect 280 61 286 65
rect 280 65 281 66
rect 282 65 283 66
rect 283 65 284 66
rect 285 65 286 66
rect 540 500 541 501
rect 542 500 543 501
rect 543 500 544 501
rect 545 500 546 501
rect 540 501 546 505
rect 540 505 541 506
rect 542 505 543 506
rect 543 505 544 506
rect 545 505 546 506
rect 400 360 401 361
rect 402 360 403 361
rect 403 360 404 361
rect 405 360 406 361
rect 400 361 406 365
rect 400 365 401 366
rect 402 365 403 366
rect 403 365 404 366
rect 405 365 406 366
rect 460 140 461 141
rect 462 140 463 141
rect 463 140 464 141
rect 465 140 466 141
rect 460 141 466 145
rect 460 145 461 146
rect 462 145 463 146
rect 463 145 464 146
rect 465 145 466 146
rect 300 180 301 181
rect 302 180 303 181
rect 303 180 304 181
rect 305 180 306 181
rect 300 181 306 185
rect 300 185 301 186
rect 302 185 303 186
rect 303 185 304 186
rect 305 185 306 186
rect 340 240 341 241
rect 342 240 343 241
rect 343 240 344 241
rect 345 240 346 241
rect 340 241 346 245
rect 340 245 341 246
rect 342 245 343 246
rect 343 245 344 246
rect 345 245 346 246
rect 200 40 201 41
rect 202 40 203 41
rect 203 40 204 41
rect 205 40 206 41
rect 200 41 206 45
rect 200 45 201 46
rect 202 45 203 46
rect 203 45 204 46
rect 205 45 206 46
rect 260 380 261 381
rect 262 380 263 381
rect 263 380 264 381
rect 265 380 266 381
rect 260 381 266 385
rect 260 385 261 386
rect 262 385 263 386
rect 263 385 264 386
rect 265 385 266 386
rect 500 560 501 561
rect 502 560 503 561
rect 503 560 504 561
rect 505 560 506 561
rect 500 561 506 565
rect 500 565 501 566
rect 502 565 503 566
rect 503 565 504 566
rect 505 565 506 566
rect 220 160 221 161
rect 222 160 223 161
rect 223 160 224 161
rect 225 160 226 161
rect 220 161 226 165
rect 220 165 221 166
rect 222 165 223 166
rect 223 165 224 166
rect 225 165 226 166
rect 280 520 281 521
rect 282 520 283 521
rect 283 520 284 521
rect 285 520 286 521
rect 280 521 286 525
rect 280 525 281 526
rect 282 525 283 526
rect 283 525 284 526
rect 285 525 286 526
rect 200 480 201 481
rect 202 480 203 481
rect 203 480 204 481
rect 205 480 206 481
rect 200 481 206 485
rect 200 485 201 486
rect 202 485 203 486
rect 203 485 204 486
rect 205 485 206 486
rect 460 60 461 61
rect 462 60 463 61
rect 463 60 464 61
rect 465 60 466 61
rect 460 61 466 65
rect 460 65 461 66
rect 462 65 463 66
rect 463 65 464 66
rect 465 65 466 66
rect 180 460 181 461
rect 182 460 183 461
rect 183 460 184 461
rect 185 460 186 461
rect 180 461 186 465
rect 180 465 181 466
rect 182 465 183 466
rect 183 465 184 466
rect 185 465 186 466
rect 320 20 321 21
rect 322 20 323 21
rect 323 20 324 21
rect 325 20 326 21
rect 320 21 326 25
rect 320 25 321 26
rect 322 25 323 26
rect 323 25 324 26
rect 325 25 326 26
rect 320 280 321 281
rect 322 280 323 281
rect 323 280 324 281
rect 325 280 326 281
rect 320 281 326 285
rect 320 285 321 286
rect 322 285 323 286
rect 323 285 324 286
rect 325 285 326 286
rect 560 260 561 261
rect 562 260 563 261
rect 563 260 564 261
rect 565 260 566 261
rect 560 261 566 265
rect 560 265 561 266
rect 562 265 563 266
rect 563 265 564 266
rect 565 265 566 266
rect 560 320 561 321
rect 562 320 563 321
rect 563 320 564 321
rect 565 320 566 321
rect 560 321 566 325
rect 560 325 561 326
rect 562 325 563 326
rect 563 325 564 326
rect 565 325 566 326
rect 660 360 661 361
rect 662 360 663 361
rect 663 360 664 361
rect 665 360 666 361
rect 660 361 666 365
rect 660 365 661 366
rect 662 365 663 366
rect 663 365 664 366
rect 665 365 666 366
rect 340 100 341 101
rect 342 100 343 101
rect 343 100 344 101
rect 345 100 346 101
rect 340 101 346 105
rect 340 105 341 106
rect 342 105 343 106
rect 343 105 344 106
rect 345 105 346 106
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect 380 140 381 141
rect 382 140 383 141
rect 383 140 384 141
rect 385 140 386 141
rect 380 141 386 145
rect 380 145 381 146
rect 382 145 383 146
rect 383 145 384 146
rect 385 145 386 146
rect 140 380 141 381
rect 142 380 143 381
rect 143 380 144 381
rect 145 380 146 381
rect 140 381 146 385
rect 140 385 141 386
rect 142 385 143 386
rect 143 385 144 386
rect 145 385 146 386
rect 320 0 321 1
rect 322 0 323 1
rect 323 0 324 1
rect 325 0 326 1
rect 320 1 326 5
rect 320 5 321 6
rect 322 5 323 6
rect 323 5 324 6
rect 325 5 326 6
rect 340 400 341 401
rect 342 400 343 401
rect 343 400 344 401
rect 345 400 346 401
rect 340 401 346 405
rect 340 405 341 406
rect 342 405 343 406
rect 343 405 344 406
rect 345 405 346 406
rect 480 400 481 401
rect 482 400 483 401
rect 483 400 484 401
rect 485 400 486 401
rect 480 401 486 405
rect 480 405 481 406
rect 482 405 483 406
rect 483 405 484 406
rect 485 405 486 406
rect 160 520 161 521
rect 162 520 163 521
rect 163 520 164 521
rect 165 520 166 521
rect 160 521 166 525
rect 160 525 161 526
rect 162 525 163 526
rect 163 525 164 526
rect 165 525 166 526
rect 280 380 281 381
rect 282 380 283 381
rect 283 380 284 381
rect 285 380 286 381
rect 280 381 286 385
rect 280 385 281 386
rect 282 385 283 386
rect 283 385 284 386
rect 285 385 286 386
rect 420 420 421 421
rect 422 420 423 421
rect 423 420 424 421
rect 425 420 426 421
rect 420 421 426 425
rect 420 425 421 426
rect 422 425 423 426
rect 423 425 424 426
rect 425 425 426 426
rect 540 540 541 541
rect 542 540 543 541
rect 543 540 544 541
rect 545 540 546 541
rect 540 541 546 545
rect 540 545 541 546
rect 542 545 543 546
rect 543 545 544 546
rect 545 545 546 546
rect 140 520 141 521
rect 142 520 143 521
rect 143 520 144 521
rect 145 520 146 521
rect 140 521 146 525
rect 140 525 141 526
rect 142 525 143 526
rect 143 525 144 526
rect 145 525 146 526
rect 460 200 461 201
rect 462 200 463 201
rect 463 200 464 201
rect 465 200 466 201
rect 460 201 466 205
rect 460 205 461 206
rect 462 205 463 206
rect 463 205 464 206
rect 465 205 466 206
rect 380 540 381 541
rect 382 540 383 541
rect 383 540 384 541
rect 385 540 386 541
rect 380 541 386 545
rect 380 545 381 546
rect 382 545 383 546
rect 383 545 384 546
rect 385 545 386 546
rect 460 180 461 181
rect 462 180 463 181
rect 463 180 464 181
rect 465 180 466 181
rect 460 181 466 185
rect 460 185 461 186
rect 462 185 463 186
rect 463 185 464 186
rect 465 185 466 186
rect 60 400 61 401
rect 62 400 63 401
rect 63 400 64 401
rect 65 400 66 401
rect 60 401 66 405
rect 60 405 61 406
rect 62 405 63 406
rect 63 405 64 406
rect 65 405 66 406
rect 240 140 241 141
rect 242 140 243 141
rect 243 140 244 141
rect 245 140 246 141
rect 240 141 246 145
rect 240 145 241 146
rect 242 145 243 146
rect 243 145 244 146
rect 245 145 246 146
rect 20 280 21 281
rect 22 280 23 281
rect 23 280 24 281
rect 25 280 26 281
rect 20 281 26 285
rect 20 285 21 286
rect 22 285 23 286
rect 23 285 24 286
rect 25 285 26 286
rect 480 600 481 601
rect 482 600 483 601
rect 483 600 484 601
rect 485 600 486 601
rect 480 601 486 605
rect 480 605 481 606
rect 482 605 483 606
rect 483 605 484 606
rect 485 605 486 606
rect 380 360 381 361
rect 382 360 383 361
rect 383 360 384 361
rect 385 360 386 361
rect 380 361 386 365
rect 380 365 381 366
rect 382 365 383 366
rect 383 365 384 366
rect 385 365 386 366
rect 240 120 241 121
rect 242 120 243 121
rect 243 120 244 121
rect 245 120 246 121
rect 240 121 246 125
rect 240 125 241 126
rect 242 125 243 126
rect 243 125 244 126
rect 245 125 246 126
rect 420 640 421 641
rect 422 640 423 641
rect 423 640 424 641
rect 425 640 426 641
rect 420 641 426 645
rect 420 645 421 646
rect 422 645 423 646
rect 423 645 424 646
rect 425 645 426 646
rect 600 160 601 161
rect 602 160 603 161
rect 603 160 604 161
rect 605 160 606 161
rect 600 161 606 165
rect 600 165 601 166
rect 602 165 603 166
rect 603 165 604 166
rect 605 165 606 166
rect 380 660 381 661
rect 382 660 383 661
rect 383 660 384 661
rect 385 660 386 661
rect 380 661 386 665
rect 380 665 381 666
rect 382 665 383 666
rect 383 665 384 666
rect 385 665 386 666
rect 280 120 281 121
rect 282 120 283 121
rect 283 120 284 121
rect 285 120 286 121
rect 280 121 286 125
rect 280 125 281 126
rect 282 125 283 126
rect 283 125 284 126
rect 285 125 286 126
rect 300 440 301 441
rect 302 440 303 441
rect 303 440 304 441
rect 305 440 306 441
rect 300 441 306 445
rect 300 445 301 446
rect 302 445 303 446
rect 303 445 304 446
rect 305 445 306 446
rect 280 540 281 541
rect 282 540 283 541
rect 283 540 284 541
rect 285 540 286 541
rect 280 541 286 545
rect 280 545 281 546
rect 282 545 283 546
rect 283 545 284 546
rect 285 545 286 546
rect 200 80 201 81
rect 202 80 203 81
rect 203 80 204 81
rect 205 80 206 81
rect 200 81 206 85
rect 200 85 201 86
rect 202 85 203 86
rect 203 85 204 86
rect 205 85 206 86
rect 20 180 21 181
rect 22 180 23 181
rect 23 180 24 181
rect 25 180 26 181
rect 20 181 26 185
rect 20 185 21 186
rect 22 185 23 186
rect 23 185 24 186
rect 25 185 26 186
rect 400 100 401 101
rect 402 100 403 101
rect 403 100 404 101
rect 405 100 406 101
rect 400 101 406 105
rect 400 105 401 106
rect 402 105 403 106
rect 403 105 404 106
rect 405 105 406 106
rect 480 640 481 641
rect 482 640 483 641
rect 483 640 484 641
rect 485 640 486 641
rect 480 641 486 645
rect 480 645 481 646
rect 482 645 483 646
rect 483 645 484 646
rect 485 645 486 646
rect 360 520 361 521
rect 362 520 363 521
rect 363 520 364 521
rect 365 520 366 521
rect 360 521 366 525
rect 360 525 361 526
rect 362 525 363 526
rect 363 525 364 526
rect 365 525 366 526
rect 80 120 81 121
rect 82 120 83 121
rect 83 120 84 121
rect 85 120 86 121
rect 80 121 86 125
rect 80 125 81 126
rect 82 125 83 126
rect 83 125 84 126
rect 85 125 86 126
rect 320 120 321 121
rect 322 120 323 121
rect 323 120 324 121
rect 325 120 326 121
rect 320 121 326 125
rect 320 125 321 126
rect 322 125 323 126
rect 323 125 324 126
rect 325 125 326 126
rect 300 200 301 201
rect 302 200 303 201
rect 303 200 304 201
rect 305 200 306 201
rect 300 201 306 205
rect 300 205 301 206
rect 302 205 303 206
rect 303 205 304 206
rect 305 205 306 206
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect 300 480 301 481
rect 302 480 303 481
rect 303 480 304 481
rect 305 480 306 481
rect 300 481 306 485
rect 300 485 301 486
rect 302 485 303 486
rect 303 485 304 486
rect 305 485 306 486
rect 40 340 41 341
rect 42 340 43 341
rect 43 340 44 341
rect 45 340 46 341
rect 40 341 46 345
rect 40 345 41 346
rect 42 345 43 346
rect 43 345 44 346
rect 45 345 46 346
rect 480 240 481 241
rect 482 240 483 241
rect 483 240 484 241
rect 485 240 486 241
rect 480 241 486 245
rect 480 245 481 246
rect 482 245 483 246
rect 483 245 484 246
rect 485 245 486 246
rect 200 260 201 261
rect 202 260 203 261
rect 203 260 204 261
rect 205 260 206 261
rect 200 261 206 265
rect 200 265 201 266
rect 202 265 203 266
rect 203 265 204 266
rect 205 265 206 266
rect 380 440 381 441
rect 382 440 383 441
rect 383 440 384 441
rect 385 440 386 441
rect 380 441 386 445
rect 380 445 381 446
rect 382 445 383 446
rect 383 445 384 446
rect 385 445 386 446
rect 280 300 281 301
rect 282 300 283 301
rect 283 300 284 301
rect 285 300 286 301
rect 280 301 286 305
rect 280 305 281 306
rect 282 305 283 306
rect 283 305 284 306
rect 285 305 286 306
rect 620 200 621 201
rect 622 200 623 201
rect 623 200 624 201
rect 625 200 626 201
rect 620 201 626 205
rect 620 205 621 206
rect 622 205 623 206
rect 623 205 624 206
rect 625 205 626 206
rect 320 480 321 481
rect 322 480 323 481
rect 323 480 324 481
rect 325 480 326 481
rect 320 481 326 485
rect 320 485 321 486
rect 322 485 323 486
rect 323 485 324 486
rect 325 485 326 486
rect 600 520 601 521
rect 602 520 603 521
rect 603 520 604 521
rect 605 520 606 521
rect 600 521 606 525
rect 600 525 601 526
rect 602 525 603 526
rect 603 525 604 526
rect 605 525 606 526
rect 120 620 121 621
rect 122 620 123 621
rect 123 620 124 621
rect 125 620 126 621
rect 120 621 126 625
rect 120 625 121 626
rect 122 625 123 626
rect 123 625 124 626
rect 125 625 126 626
rect 400 200 401 201
rect 402 200 403 201
rect 403 200 404 201
rect 405 200 406 201
rect 400 201 406 205
rect 400 205 401 206
rect 402 205 403 206
rect 403 205 404 206
rect 405 205 406 206
rect 20 400 21 401
rect 22 400 23 401
rect 23 400 24 401
rect 25 400 26 401
rect 20 401 26 405
rect 20 405 21 406
rect 22 405 23 406
rect 23 405 24 406
rect 25 405 26 406
rect 280 0 281 1
rect 282 0 283 1
rect 283 0 284 1
rect 285 0 286 1
rect 280 1 286 5
rect 280 5 281 6
rect 282 5 283 6
rect 283 5 284 6
rect 285 5 286 6
rect 280 400 281 401
rect 282 400 283 401
rect 283 400 284 401
rect 285 400 286 401
rect 280 401 286 405
rect 280 405 281 406
rect 282 405 283 406
rect 283 405 284 406
rect 285 405 286 406
rect 460 240 461 241
rect 462 240 463 241
rect 463 240 464 241
rect 465 240 466 241
rect 460 241 466 245
rect 460 245 461 246
rect 462 245 463 246
rect 463 245 464 246
rect 465 245 466 246
rect 300 280 301 281
rect 302 280 303 281
rect 303 280 304 281
rect 305 280 306 281
rect 300 281 306 285
rect 300 285 301 286
rect 302 285 303 286
rect 303 285 304 286
rect 305 285 306 286
rect 440 600 441 601
rect 442 600 443 601
rect 443 600 444 601
rect 445 600 446 601
rect 440 601 446 605
rect 440 605 441 606
rect 442 605 443 606
rect 443 605 444 606
rect 445 605 446 606
rect 120 420 121 421
rect 122 420 123 421
rect 123 420 124 421
rect 125 420 126 421
rect 120 421 126 425
rect 120 425 121 426
rect 122 425 123 426
rect 123 425 124 426
rect 125 425 126 426
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect 100 540 101 541
rect 102 540 103 541
rect 103 540 104 541
rect 105 540 106 541
rect 100 541 106 545
rect 100 545 101 546
rect 102 545 103 546
rect 103 545 104 546
rect 105 545 106 546
rect 340 80 341 81
rect 342 80 343 81
rect 343 80 344 81
rect 345 80 346 81
rect 340 81 346 85
rect 340 85 341 86
rect 342 85 343 86
rect 343 85 344 86
rect 345 85 346 86
rect 220 440 221 441
rect 222 440 223 441
rect 223 440 224 441
rect 225 440 226 441
rect 220 441 226 445
rect 220 445 221 446
rect 222 445 223 446
rect 223 445 224 446
rect 225 445 226 446
rect 340 180 341 181
rect 342 180 343 181
rect 343 180 344 181
rect 345 180 346 181
rect 340 181 346 185
rect 340 185 341 186
rect 342 185 343 186
rect 343 185 344 186
rect 345 185 346 186
rect 360 320 361 321
rect 362 320 363 321
rect 363 320 364 321
rect 365 320 366 321
rect 360 321 366 325
rect 360 325 361 326
rect 362 325 363 326
rect 363 325 364 326
rect 365 325 366 326
rect 40 240 41 241
rect 42 240 43 241
rect 43 240 44 241
rect 45 240 46 241
rect 40 241 46 245
rect 40 245 41 246
rect 42 245 43 246
rect 43 245 44 246
rect 45 245 46 246
rect 180 660 181 661
rect 182 660 183 661
rect 183 660 184 661
rect 185 660 186 661
rect 180 661 186 665
rect 180 665 181 666
rect 182 665 183 666
rect 183 665 184 666
rect 185 665 186 666
rect 520 40 521 41
rect 522 40 523 41
rect 523 40 524 41
rect 525 40 526 41
rect 520 41 526 45
rect 520 45 521 46
rect 522 45 523 46
rect 523 45 524 46
rect 525 45 526 46
rect 240 300 241 301
rect 242 300 243 301
rect 243 300 244 301
rect 245 300 246 301
rect 240 301 246 305
rect 240 305 241 306
rect 242 305 243 306
rect 243 305 244 306
rect 245 305 246 306
rect 360 160 361 161
rect 362 160 363 161
rect 363 160 364 161
rect 365 160 366 161
rect 360 161 366 165
rect 360 165 361 166
rect 362 165 363 166
rect 363 165 364 166
rect 365 165 366 166
rect 400 520 401 521
rect 402 520 403 521
rect 403 520 404 521
rect 405 520 406 521
rect 400 521 406 525
rect 400 525 401 526
rect 402 525 403 526
rect 403 525 404 526
rect 405 525 406 526
rect 340 640 341 641
rect 342 640 343 641
rect 343 640 344 641
rect 345 640 346 641
rect 340 641 346 645
rect 340 645 341 646
rect 342 645 343 646
rect 343 645 344 646
rect 345 645 346 646
rect 200 160 201 161
rect 202 160 203 161
rect 203 160 204 161
rect 205 160 206 161
rect 200 161 206 165
rect 200 165 201 166
rect 202 165 203 166
rect 203 165 204 166
rect 205 165 206 166
rect 20 100 21 101
rect 22 100 23 101
rect 23 100 24 101
rect 25 100 26 101
rect 20 101 26 105
rect 20 105 21 106
rect 22 105 23 106
rect 23 105 24 106
rect 25 105 26 106
rect 340 480 341 481
rect 342 480 343 481
rect 343 480 344 481
rect 345 480 346 481
rect 340 481 346 485
rect 340 485 341 486
rect 342 485 343 486
rect 343 485 344 486
rect 345 485 346 486
rect 160 260 161 261
rect 162 260 163 261
rect 163 260 164 261
rect 165 260 166 261
rect 160 261 166 265
rect 160 265 161 266
rect 162 265 163 266
rect 163 265 164 266
rect 165 265 166 266
rect 500 140 501 141
rect 502 140 503 141
rect 503 140 504 141
rect 505 140 506 141
rect 500 141 506 145
rect 500 145 501 146
rect 502 145 503 146
rect 503 145 504 146
rect 505 145 506 146
rect 400 40 401 41
rect 402 40 403 41
rect 403 40 404 41
rect 405 40 406 41
rect 400 41 406 45
rect 400 45 401 46
rect 402 45 403 46
rect 403 45 404 46
rect 405 45 406 46
rect 240 540 241 541
rect 242 540 243 541
rect 243 540 244 541
rect 245 540 246 541
rect 240 541 246 545
rect 240 545 241 546
rect 242 545 243 546
rect 243 545 244 546
rect 245 545 246 546
rect 520 540 521 541
rect 522 540 523 541
rect 523 540 524 541
rect 525 540 526 541
rect 520 541 526 545
rect 520 545 521 546
rect 522 545 523 546
rect 523 545 524 546
rect 525 545 526 546
rect 340 320 341 321
rect 342 320 343 321
rect 343 320 344 321
rect 345 320 346 321
rect 340 321 346 325
rect 340 325 341 326
rect 342 325 343 326
rect 343 325 344 326
rect 345 325 346 326
rect 380 460 381 461
rect 382 460 383 461
rect 383 460 384 461
rect 385 460 386 461
rect 380 461 386 465
rect 380 465 381 466
rect 382 465 383 466
rect 383 465 384 466
rect 385 465 386 466
rect 100 220 101 221
rect 102 220 103 221
rect 103 220 104 221
rect 105 220 106 221
rect 100 221 106 225
rect 100 225 101 226
rect 102 225 103 226
rect 103 225 104 226
rect 105 225 106 226
rect 600 180 601 181
rect 602 180 603 181
rect 603 180 604 181
rect 605 180 606 181
rect 600 181 606 185
rect 600 185 601 186
rect 602 185 603 186
rect 603 185 604 186
rect 605 185 606 186
rect 460 340 461 341
rect 462 340 463 341
rect 463 340 464 341
rect 465 340 466 341
rect 460 341 466 345
rect 460 345 461 346
rect 462 345 463 346
rect 463 345 464 346
rect 465 345 466 346
rect 80 160 81 161
rect 82 160 83 161
rect 83 160 84 161
rect 85 160 86 161
rect 80 161 86 165
rect 80 165 81 166
rect 82 165 83 166
rect 83 165 84 166
rect 85 165 86 166
rect 520 200 521 201
rect 522 200 523 201
rect 523 200 524 201
rect 525 200 526 201
rect 520 201 526 205
rect 520 205 521 206
rect 522 205 523 206
rect 523 205 524 206
rect 525 205 526 206
rect 200 360 201 361
rect 202 360 203 361
rect 203 360 204 361
rect 205 360 206 361
rect 200 361 206 365
rect 200 365 201 366
rect 202 365 203 366
rect 203 365 204 366
rect 205 365 206 366
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect 120 140 121 141
rect 122 140 123 141
rect 123 140 124 141
rect 125 140 126 141
rect 120 141 126 145
rect 120 145 121 146
rect 122 145 123 146
rect 123 145 124 146
rect 125 145 126 146
rect 160 420 161 421
rect 162 420 163 421
rect 163 420 164 421
rect 165 420 166 421
rect 160 421 166 425
rect 160 425 161 426
rect 162 425 163 426
rect 163 425 164 426
rect 165 425 166 426
rect 320 400 321 401
rect 322 400 323 401
rect 323 400 324 401
rect 325 400 326 401
rect 320 401 326 405
rect 320 405 321 406
rect 322 405 323 406
rect 323 405 324 406
rect 325 405 326 406
rect 460 520 461 521
rect 462 520 463 521
rect 463 520 464 521
rect 465 520 466 521
rect 460 521 466 525
rect 460 525 461 526
rect 462 525 463 526
rect 463 525 464 526
rect 465 525 466 526
rect 360 380 361 381
rect 362 380 363 381
rect 363 380 364 381
rect 365 380 366 381
rect 360 381 366 385
rect 360 385 361 386
rect 362 385 363 386
rect 363 385 364 386
rect 365 385 366 386
rect 260 440 261 441
rect 262 440 263 441
rect 263 440 264 441
rect 265 440 266 441
rect 260 441 266 445
rect 260 445 261 446
rect 262 445 263 446
rect 263 445 264 446
rect 265 445 266 446
rect 280 440 281 441
rect 282 440 283 441
rect 283 440 284 441
rect 285 440 286 441
rect 280 441 286 445
rect 280 445 281 446
rect 282 445 283 446
rect 283 445 284 446
rect 285 445 286 446
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect 500 380 501 381
rect 502 380 503 381
rect 503 380 504 381
rect 505 380 506 381
rect 500 381 506 385
rect 500 385 501 386
rect 502 385 503 386
rect 503 385 504 386
rect 505 385 506 386
rect 500 340 501 341
rect 502 340 503 341
rect 503 340 504 341
rect 505 340 506 341
rect 500 341 506 345
rect 500 345 501 346
rect 502 345 503 346
rect 503 345 504 346
rect 505 345 506 346
rect 340 540 341 541
rect 342 540 343 541
rect 343 540 344 541
rect 345 540 346 541
rect 340 541 346 545
rect 340 545 341 546
rect 342 545 343 546
rect 343 545 344 546
rect 345 545 346 546
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect 540 380 541 381
rect 542 380 543 381
rect 543 380 544 381
rect 545 380 546 381
rect 540 381 546 385
rect 540 385 541 386
rect 542 385 543 386
rect 543 385 544 386
rect 545 385 546 386
rect 260 260 261 261
rect 262 260 263 261
rect 263 260 264 261
rect 265 260 266 261
rect 260 261 266 265
rect 260 265 261 266
rect 262 265 263 266
rect 263 265 264 266
rect 265 265 266 266
rect 440 220 441 221
rect 442 220 443 221
rect 443 220 444 221
rect 445 220 446 221
rect 440 221 446 225
rect 440 225 441 226
rect 442 225 443 226
rect 443 225 444 226
rect 445 225 446 226
rect 160 240 161 241
rect 162 240 163 241
rect 163 240 164 241
rect 165 240 166 241
rect 160 241 166 245
rect 160 245 161 246
rect 162 245 163 246
rect 163 245 164 246
rect 165 245 166 246
rect 480 540 481 541
rect 482 540 483 541
rect 483 540 484 541
rect 485 540 486 541
rect 480 541 486 545
rect 480 545 481 546
rect 482 545 483 546
rect 483 545 484 546
rect 485 545 486 546
rect 380 560 381 561
rect 382 560 383 561
rect 383 560 384 561
rect 385 560 386 561
rect 380 561 386 565
rect 380 565 381 566
rect 382 565 383 566
rect 383 565 384 566
rect 385 565 386 566
rect 440 400 441 401
rect 442 400 443 401
rect 443 400 444 401
rect 445 400 446 401
rect 440 401 446 405
rect 440 405 441 406
rect 442 405 443 406
rect 443 405 444 406
rect 445 405 446 406
rect 620 180 621 181
rect 622 180 623 181
rect 623 180 624 181
rect 625 180 626 181
rect 620 181 626 185
rect 620 185 621 186
rect 622 185 623 186
rect 623 185 624 186
rect 625 185 626 186
rect 300 300 301 301
rect 302 300 303 301
rect 303 300 304 301
rect 305 300 306 301
rect 300 301 306 305
rect 300 305 301 306
rect 302 305 303 306
rect 303 305 304 306
rect 305 305 306 306
rect 540 600 541 601
rect 542 600 543 601
rect 543 600 544 601
rect 545 600 546 601
rect 540 601 546 605
rect 540 605 541 606
rect 542 605 543 606
rect 543 605 544 606
rect 545 605 546 606
rect 20 240 21 241
rect 22 240 23 241
rect 23 240 24 241
rect 25 240 26 241
rect 20 241 26 245
rect 20 245 21 246
rect 22 245 23 246
rect 23 245 24 246
rect 25 245 26 246
rect 320 540 321 541
rect 322 540 323 541
rect 323 540 324 541
rect 325 540 326 541
rect 320 541 326 545
rect 320 545 321 546
rect 322 545 323 546
rect 323 545 324 546
rect 325 545 326 546
rect 360 660 361 661
rect 362 660 363 661
rect 363 660 364 661
rect 365 660 366 661
rect 360 661 366 665
rect 360 665 361 666
rect 362 665 363 666
rect 363 665 364 666
rect 365 665 366 666
rect 280 340 281 341
rect 282 340 283 341
rect 283 340 284 341
rect 285 340 286 341
rect 280 341 286 345
rect 280 345 281 346
rect 282 345 283 346
rect 283 345 284 346
rect 285 345 286 346
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect 440 460 441 461
rect 442 460 443 461
rect 443 460 444 461
rect 445 460 446 461
rect 440 461 446 465
rect 440 465 441 466
rect 442 465 443 466
rect 443 465 444 466
rect 445 465 446 466
rect 260 140 261 141
rect 262 140 263 141
rect 263 140 264 141
rect 265 140 266 141
rect 260 141 266 145
rect 260 145 261 146
rect 262 145 263 146
rect 263 145 264 146
rect 265 145 266 146
rect 580 240 581 241
rect 582 240 583 241
rect 583 240 584 241
rect 585 240 586 241
rect 580 241 586 245
rect 580 245 581 246
rect 582 245 583 246
rect 583 245 584 246
rect 585 245 586 246
rect 220 60 221 61
rect 222 60 223 61
rect 223 60 224 61
rect 225 60 226 61
rect 220 61 226 65
rect 220 65 221 66
rect 222 65 223 66
rect 223 65 224 66
rect 225 65 226 66
rect 400 540 401 541
rect 402 540 403 541
rect 403 540 404 541
rect 405 540 406 541
rect 400 541 406 545
rect 400 545 401 546
rect 402 545 403 546
rect 403 545 404 546
rect 405 545 406 546
rect 280 420 281 421
rect 282 420 283 421
rect 283 420 284 421
rect 285 420 286 421
rect 280 421 286 425
rect 280 425 281 426
rect 282 425 283 426
rect 283 425 284 426
rect 285 425 286 426
rect 320 500 321 501
rect 322 500 323 501
rect 323 500 324 501
rect 325 500 326 501
rect 320 501 326 505
rect 320 505 321 506
rect 322 505 323 506
rect 323 505 324 506
rect 325 505 326 506
rect 320 460 321 461
rect 322 460 323 461
rect 323 460 324 461
rect 325 460 326 461
rect 320 461 326 465
rect 320 465 321 466
rect 322 465 323 466
rect 323 465 324 466
rect 325 465 326 466
rect 0 260 1 261
rect 2 260 3 261
rect 3 260 4 261
rect 5 260 6 261
rect 0 261 6 265
rect 0 265 1 266
rect 2 265 3 266
rect 3 265 4 266
rect 5 265 6 266
rect 240 460 241 461
rect 242 460 243 461
rect 243 460 244 461
rect 245 460 246 461
rect 240 461 246 465
rect 240 465 241 466
rect 242 465 243 466
rect 243 465 244 466
rect 245 465 246 466
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect 140 120 141 121
rect 142 120 143 121
rect 143 120 144 121
rect 145 120 146 121
rect 140 121 146 125
rect 140 125 141 126
rect 142 125 143 126
rect 143 125 144 126
rect 145 125 146 126
rect 560 180 561 181
rect 562 180 563 181
rect 563 180 564 181
rect 565 180 566 181
rect 560 181 566 185
rect 560 185 561 186
rect 562 185 563 186
rect 563 185 564 186
rect 565 185 566 186
rect 60 160 61 161
rect 62 160 63 161
rect 63 160 64 161
rect 65 160 66 161
rect 60 161 66 165
rect 60 165 61 166
rect 62 165 63 166
rect 63 165 64 166
rect 65 165 66 166
rect 520 140 521 141
rect 522 140 523 141
rect 523 140 524 141
rect 525 140 526 141
rect 520 141 526 145
rect 520 145 521 146
rect 522 145 523 146
rect 523 145 524 146
rect 525 145 526 146
rect 260 340 261 341
rect 262 340 263 341
rect 263 340 264 341
rect 265 340 266 341
rect 260 341 266 345
rect 260 345 261 346
rect 262 345 263 346
rect 263 345 264 346
rect 265 345 266 346
rect 320 220 321 221
rect 322 220 323 221
rect 323 220 324 221
rect 325 220 326 221
rect 320 221 326 225
rect 320 225 321 226
rect 322 225 323 226
rect 323 225 324 226
rect 325 225 326 226
rect 440 440 441 441
rect 442 440 443 441
rect 443 440 444 441
rect 445 440 446 441
rect 440 441 446 445
rect 440 445 441 446
rect 442 445 443 446
rect 443 445 444 446
rect 445 445 446 446
rect 200 640 201 641
rect 202 640 203 641
rect 203 640 204 641
rect 205 640 206 641
rect 200 641 206 645
rect 200 645 201 646
rect 202 645 203 646
rect 203 645 204 646
rect 205 645 206 646
rect 360 500 361 501
rect 362 500 363 501
rect 363 500 364 501
rect 365 500 366 501
rect 360 501 366 505
rect 360 505 361 506
rect 362 505 363 506
rect 363 505 364 506
rect 365 505 366 506
rect 20 500 21 501
rect 22 500 23 501
rect 23 500 24 501
rect 25 500 26 501
rect 20 501 26 505
rect 20 505 21 506
rect 22 505 23 506
rect 23 505 24 506
rect 25 505 26 506
rect 380 60 381 61
rect 382 60 383 61
rect 383 60 384 61
rect 385 60 386 61
rect 380 61 386 65
rect 380 65 381 66
rect 382 65 383 66
rect 383 65 384 66
rect 385 65 386 66
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect 340 220 341 221
rect 342 220 343 221
rect 343 220 344 221
rect 345 220 346 221
rect 340 221 346 225
rect 340 225 341 226
rect 342 225 343 226
rect 343 225 344 226
rect 345 225 346 226
rect 460 380 461 381
rect 462 380 463 381
rect 463 380 464 381
rect 465 380 466 381
rect 460 381 466 385
rect 460 385 461 386
rect 462 385 463 386
rect 463 385 464 386
rect 465 385 466 386
rect 660 280 661 281
rect 662 280 663 281
rect 663 280 664 281
rect 665 280 666 281
rect 660 281 666 285
rect 660 285 661 286
rect 662 285 663 286
rect 663 285 664 286
rect 665 285 666 286
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect 40 260 41 261
rect 42 260 43 261
rect 43 260 44 261
rect 45 260 46 261
rect 40 261 46 265
rect 40 265 41 266
rect 42 265 43 266
rect 43 265 44 266
rect 45 265 46 266
rect 240 480 241 481
rect 242 480 243 481
rect 243 480 244 481
rect 245 480 246 481
rect 240 481 246 485
rect 240 485 241 486
rect 242 485 243 486
rect 243 485 244 486
rect 245 485 246 486
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect 660 340 661 341
rect 662 340 663 341
rect 663 340 664 341
rect 665 340 666 341
rect 660 341 666 345
rect 660 345 661 346
rect 662 345 663 346
rect 663 345 664 346
rect 665 345 666 346
rect 140 440 141 441
rect 142 440 143 441
rect 143 440 144 441
rect 145 440 146 441
rect 140 441 146 445
rect 140 445 141 446
rect 142 445 143 446
rect 143 445 144 446
rect 145 445 146 446
rect 520 100 521 101
rect 522 100 523 101
rect 523 100 524 101
rect 525 100 526 101
rect 520 101 526 105
rect 520 105 521 106
rect 522 105 523 106
rect 523 105 524 106
rect 525 105 526 106
rect 620 400 621 401
rect 622 400 623 401
rect 623 400 624 401
rect 625 400 626 401
rect 620 401 626 405
rect 620 405 621 406
rect 622 405 623 406
rect 623 405 624 406
rect 625 405 626 406
rect 280 320 281 321
rect 282 320 283 321
rect 283 320 284 321
rect 285 320 286 321
rect 280 321 286 325
rect 280 325 281 326
rect 282 325 283 326
rect 283 325 284 326
rect 285 325 286 326
rect 60 120 61 121
rect 62 120 63 121
rect 63 120 64 121
rect 65 120 66 121
rect 60 121 66 125
rect 60 125 61 126
rect 62 125 63 126
rect 63 125 64 126
rect 65 125 66 126
rect 340 120 341 121
rect 342 120 343 121
rect 343 120 344 121
rect 345 120 346 121
rect 340 121 346 125
rect 340 125 341 126
rect 342 125 343 126
rect 343 125 344 126
rect 345 125 346 126
rect 440 340 441 341
rect 442 340 443 341
rect 443 340 444 341
rect 445 340 446 341
rect 440 341 446 345
rect 440 345 441 346
rect 442 345 443 346
rect 443 345 444 346
rect 445 345 446 346
rect 520 360 521 361
rect 522 360 523 361
rect 523 360 524 361
rect 525 360 526 361
rect 520 361 526 365
rect 520 365 521 366
rect 522 365 523 366
rect 523 365 524 366
rect 525 365 526 366
rect 320 380 321 381
rect 322 380 323 381
rect 323 380 324 381
rect 325 380 326 381
rect 320 381 326 385
rect 320 385 321 386
rect 322 385 323 386
rect 323 385 324 386
rect 325 385 326 386
rect 600 400 601 401
rect 602 400 603 401
rect 603 400 604 401
rect 605 400 606 401
rect 600 401 606 405
rect 600 405 601 406
rect 602 405 603 406
rect 603 405 604 406
rect 605 405 606 406
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect 600 260 601 261
rect 602 260 603 261
rect 603 260 604 261
rect 605 260 606 261
rect 600 261 606 265
rect 600 265 601 266
rect 602 265 603 266
rect 603 265 604 266
rect 605 265 606 266
rect 220 40 221 41
rect 222 40 223 41
rect 223 40 224 41
rect 225 40 226 41
rect 220 41 226 45
rect 220 45 221 46
rect 222 45 223 46
rect 223 45 224 46
rect 225 45 226 46
rect 120 120 121 121
rect 122 120 123 121
rect 123 120 124 121
rect 125 120 126 121
rect 120 121 126 125
rect 120 125 121 126
rect 122 125 123 126
rect 123 125 124 126
rect 125 125 126 126
rect 500 500 501 501
rect 502 500 503 501
rect 503 500 504 501
rect 505 500 506 501
rect 500 501 506 505
rect 500 505 501 506
rect 502 505 503 506
rect 503 505 504 506
rect 505 505 506 506
rect 140 500 141 501
rect 142 500 143 501
rect 143 500 144 501
rect 145 500 146 501
rect 140 501 146 505
rect 140 505 141 506
rect 142 505 143 506
rect 143 505 144 506
rect 145 505 146 506
rect 440 660 441 661
rect 442 660 443 661
rect 443 660 444 661
rect 445 660 446 661
rect 440 661 446 665
rect 440 665 441 666
rect 442 665 443 666
rect 443 665 444 666
rect 445 665 446 666
rect 400 340 401 341
rect 402 340 403 341
rect 403 340 404 341
rect 405 340 406 341
rect 400 341 406 345
rect 400 345 401 346
rect 402 345 403 346
rect 403 345 404 346
rect 405 345 406 346
rect 400 220 401 221
rect 402 220 403 221
rect 403 220 404 221
rect 405 220 406 221
rect 400 221 406 225
rect 400 225 401 226
rect 402 225 403 226
rect 403 225 404 226
rect 405 225 406 226
rect 120 320 121 321
rect 122 320 123 321
rect 123 320 124 321
rect 125 320 126 321
rect 120 321 126 325
rect 120 325 121 326
rect 122 325 123 326
rect 123 325 124 326
rect 125 325 126 326
rect 420 280 421 281
rect 422 280 423 281
rect 423 280 424 281
rect 425 280 426 281
rect 420 281 426 285
rect 420 285 421 286
rect 422 285 423 286
rect 423 285 424 286
rect 425 285 426 286
rect 540 220 541 221
rect 542 220 543 221
rect 543 220 544 221
rect 545 220 546 221
rect 540 221 546 225
rect 540 225 541 226
rect 542 225 543 226
rect 543 225 544 226
rect 545 225 546 226
rect 220 180 221 181
rect 222 180 223 181
rect 223 180 224 181
rect 225 180 226 181
rect 220 181 226 185
rect 220 185 221 186
rect 222 185 223 186
rect 223 185 224 186
rect 225 185 226 186
rect 280 20 281 21
rect 282 20 283 21
rect 283 20 284 21
rect 285 20 286 21
rect 280 21 286 25
rect 280 25 281 26
rect 282 25 283 26
rect 283 25 284 26
rect 285 25 286 26
rect 420 600 421 601
rect 422 600 423 601
rect 423 600 424 601
rect 425 600 426 601
rect 420 601 426 605
rect 420 605 421 606
rect 422 605 423 606
rect 423 605 424 606
rect 425 605 426 606
rect 180 120 181 121
rect 182 120 183 121
rect 183 120 184 121
rect 185 120 186 121
rect 180 121 186 125
rect 180 125 181 126
rect 182 125 183 126
rect 183 125 184 126
rect 185 125 186 126
rect 460 500 461 501
rect 462 500 463 501
rect 463 500 464 501
rect 465 500 466 501
rect 460 501 466 505
rect 460 505 461 506
rect 462 505 463 506
rect 463 505 464 506
rect 465 505 466 506
rect 240 380 241 381
rect 242 380 243 381
rect 243 380 244 381
rect 245 380 246 381
rect 240 381 246 385
rect 240 385 241 386
rect 242 385 243 386
rect 243 385 244 386
rect 245 385 246 386
rect 240 220 241 221
rect 242 220 243 221
rect 243 220 244 221
rect 245 220 246 221
rect 240 221 246 225
rect 240 225 241 226
rect 242 225 243 226
rect 243 225 244 226
rect 245 225 246 226
rect 300 340 301 341
rect 302 340 303 341
rect 303 340 304 341
rect 305 340 306 341
rect 300 341 306 345
rect 300 345 301 346
rect 302 345 303 346
rect 303 345 304 346
rect 305 345 306 346
rect 460 260 461 261
rect 462 260 463 261
rect 463 260 464 261
rect 465 260 466 261
rect 460 261 466 265
rect 460 265 461 266
rect 462 265 463 266
rect 463 265 464 266
rect 465 265 466 266
rect 120 440 121 441
rect 122 440 123 441
rect 123 440 124 441
rect 125 440 126 441
rect 120 441 126 445
rect 120 445 121 446
rect 122 445 123 446
rect 123 445 124 446
rect 125 445 126 446
rect 180 540 181 541
rect 182 540 183 541
rect 183 540 184 541
rect 185 540 186 541
rect 180 541 186 545
rect 180 545 181 546
rect 182 545 183 546
rect 183 545 184 546
rect 185 545 186 546
rect 460 80 461 81
rect 462 80 463 81
rect 463 80 464 81
rect 465 80 466 81
rect 460 81 466 85
rect 460 85 461 86
rect 462 85 463 86
rect 463 85 464 86
rect 465 85 466 86
rect 580 300 581 301
rect 582 300 583 301
rect 583 300 584 301
rect 585 300 586 301
rect 580 301 586 305
rect 580 305 581 306
rect 582 305 583 306
rect 583 305 584 306
rect 585 305 586 306
rect 460 420 461 421
rect 462 420 463 421
rect 463 420 464 421
rect 465 420 466 421
rect 460 421 466 425
rect 460 425 461 426
rect 462 425 463 426
rect 463 425 464 426
rect 465 425 466 426
rect 120 340 121 341
rect 122 340 123 341
rect 123 340 124 341
rect 125 340 126 341
rect 120 341 126 345
rect 120 345 121 346
rect 122 345 123 346
rect 123 345 124 346
rect 125 345 126 346
rect 220 320 221 321
rect 222 320 223 321
rect 223 320 224 321
rect 225 320 226 321
rect 220 321 226 325
rect 220 325 221 326
rect 222 325 223 326
rect 223 325 224 326
rect 225 325 226 326
rect 420 80 421 81
rect 422 80 423 81
rect 423 80 424 81
rect 425 80 426 81
rect 420 81 426 85
rect 420 85 421 86
rect 422 85 423 86
rect 423 85 424 86
rect 425 85 426 86
rect 60 560 61 561
rect 62 560 63 561
rect 63 560 64 561
rect 65 560 66 561
rect 60 561 66 565
rect 60 565 61 566
rect 62 565 63 566
rect 63 565 64 566
rect 65 565 66 566
rect 420 220 421 221
rect 422 220 423 221
rect 423 220 424 221
rect 425 220 426 221
rect 420 221 426 225
rect 420 225 421 226
rect 422 225 423 226
rect 423 225 424 226
rect 425 225 426 226
rect 320 520 321 521
rect 322 520 323 521
rect 323 520 324 521
rect 325 520 326 521
rect 320 521 326 525
rect 320 525 321 526
rect 322 525 323 526
rect 323 525 324 526
rect 325 525 326 526
rect 400 140 401 141
rect 402 140 403 141
rect 403 140 404 141
rect 405 140 406 141
rect 400 141 406 145
rect 400 145 401 146
rect 402 145 403 146
rect 403 145 404 146
rect 405 145 406 146
rect 400 120 401 121
rect 402 120 403 121
rect 403 120 404 121
rect 405 120 406 121
rect 400 121 406 125
rect 400 125 401 126
rect 402 125 403 126
rect 403 125 404 126
rect 405 125 406 126
rect 380 480 381 481
rect 382 480 383 481
rect 383 480 384 481
rect 385 480 386 481
rect 380 481 386 485
rect 380 485 381 486
rect 382 485 383 486
rect 383 485 384 486
rect 385 485 386 486
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect 120 100 121 101
rect 122 100 123 101
rect 123 100 124 101
rect 125 100 126 101
rect 120 101 126 105
rect 120 105 121 106
rect 122 105 123 106
rect 123 105 124 106
rect 125 105 126 106
rect 500 100 501 101
rect 502 100 503 101
rect 503 100 504 101
rect 505 100 506 101
rect 500 101 506 105
rect 500 105 501 106
rect 502 105 503 106
rect 503 105 504 106
rect 505 105 506 106
rect 300 380 301 381
rect 302 380 303 381
rect 303 380 304 381
rect 305 380 306 381
rect 300 381 306 385
rect 300 385 301 386
rect 302 385 303 386
rect 303 385 304 386
rect 305 385 306 386
rect 80 440 81 441
rect 82 440 83 441
rect 83 440 84 441
rect 85 440 86 441
rect 80 441 86 445
rect 80 445 81 446
rect 82 445 83 446
rect 83 445 84 446
rect 85 445 86 446
rect 380 600 381 601
rect 382 600 383 601
rect 383 600 384 601
rect 385 600 386 601
rect 380 601 386 605
rect 380 605 381 606
rect 382 605 383 606
rect 383 605 384 606
rect 385 605 386 606
rect 200 0 201 1
rect 202 0 203 1
rect 203 0 204 1
rect 205 0 206 1
rect 200 1 206 5
rect 200 5 201 6
rect 202 5 203 6
rect 203 5 204 6
rect 205 5 206 6
rect 480 340 481 341
rect 482 340 483 341
rect 483 340 484 341
rect 485 340 486 341
rect 480 341 486 345
rect 480 345 481 346
rect 482 345 483 346
rect 483 345 484 346
rect 485 345 486 346
rect 220 100 221 101
rect 222 100 223 101
rect 223 100 224 101
rect 225 100 226 101
rect 220 101 226 105
rect 220 105 221 106
rect 222 105 223 106
rect 223 105 224 106
rect 225 105 226 106
rect 160 160 161 161
rect 162 160 163 161
rect 163 160 164 161
rect 165 160 166 161
rect 160 161 166 165
rect 160 165 161 166
rect 162 165 163 166
rect 163 165 164 166
rect 165 165 166 166
rect 140 260 141 261
rect 142 260 143 261
rect 143 260 144 261
rect 145 260 146 261
rect 140 261 146 265
rect 140 265 141 266
rect 142 265 143 266
rect 143 265 144 266
rect 145 265 146 266
rect 100 500 101 501
rect 102 500 103 501
rect 103 500 104 501
rect 105 500 106 501
rect 100 501 106 505
rect 100 505 101 506
rect 102 505 103 506
rect 103 505 104 506
rect 105 505 106 506
rect 160 440 161 441
rect 162 440 163 441
rect 163 440 164 441
rect 165 440 166 441
rect 160 441 166 445
rect 160 445 161 446
rect 162 445 163 446
rect 163 445 164 446
rect 165 445 166 446
rect 520 580 521 581
rect 522 580 523 581
rect 523 580 524 581
rect 525 580 526 581
rect 520 581 526 585
rect 520 585 521 586
rect 522 585 523 586
rect 523 585 524 586
rect 525 585 526 586
rect 300 540 301 541
rect 302 540 303 541
rect 303 540 304 541
rect 305 540 306 541
rect 300 541 306 545
rect 300 545 301 546
rect 302 545 303 546
rect 303 545 304 546
rect 305 545 306 546
rect 380 580 381 581
rect 382 580 383 581
rect 383 580 384 581
rect 385 580 386 581
rect 380 581 386 585
rect 380 585 381 586
rect 382 585 383 586
rect 383 585 384 586
rect 385 585 386 586
rect 360 180 361 181
rect 362 180 363 181
rect 363 180 364 181
rect 365 180 366 181
rect 360 181 366 185
rect 360 185 361 186
rect 362 185 363 186
rect 363 185 364 186
rect 365 185 366 186
rect 20 220 21 221
rect 22 220 23 221
rect 23 220 24 221
rect 25 220 26 221
rect 20 221 26 225
rect 20 225 21 226
rect 22 225 23 226
rect 23 225 24 226
rect 25 225 26 226
rect 660 320 661 321
rect 662 320 663 321
rect 663 320 664 321
rect 665 320 666 321
rect 660 321 666 325
rect 660 325 661 326
rect 662 325 663 326
rect 663 325 664 326
rect 665 325 666 326
rect 320 80 321 81
rect 322 80 323 81
rect 323 80 324 81
rect 325 80 326 81
rect 320 81 326 85
rect 320 85 321 86
rect 322 85 323 86
rect 323 85 324 86
rect 325 85 326 86
rect 320 60 321 61
rect 322 60 323 61
rect 323 60 324 61
rect 325 60 326 61
rect 320 61 326 65
rect 320 65 321 66
rect 322 65 323 66
rect 323 65 324 66
rect 325 65 326 66
rect 260 580 261 581
rect 262 580 263 581
rect 263 580 264 581
rect 265 580 266 581
rect 260 581 266 585
rect 260 585 261 586
rect 262 585 263 586
rect 263 585 264 586
rect 265 585 266 586
rect 260 60 261 61
rect 262 60 263 61
rect 263 60 264 61
rect 265 60 266 61
rect 260 61 266 65
rect 260 65 261 66
rect 262 65 263 66
rect 263 65 264 66
rect 265 65 266 66
rect 220 500 221 501
rect 222 500 223 501
rect 223 500 224 501
rect 225 500 226 501
rect 220 501 226 505
rect 220 505 221 506
rect 222 505 223 506
rect 223 505 224 506
rect 225 505 226 506
rect 460 20 461 21
rect 462 20 463 21
rect 463 20 464 21
rect 465 20 466 21
rect 460 21 466 25
rect 460 25 461 26
rect 462 25 463 26
rect 463 25 464 26
rect 465 25 466 26
rect 100 400 101 401
rect 102 400 103 401
rect 103 400 104 401
rect 105 400 106 401
rect 100 401 106 405
rect 100 405 101 406
rect 102 405 103 406
rect 103 405 104 406
rect 105 405 106 406
rect 380 20 381 21
rect 382 20 383 21
rect 383 20 384 21
rect 385 20 386 21
rect 380 21 386 25
rect 380 25 381 26
rect 382 25 383 26
rect 383 25 384 26
rect 385 25 386 26
rect 260 120 261 121
rect 262 120 263 121
rect 263 120 264 121
rect 265 120 266 121
rect 260 121 266 125
rect 260 125 261 126
rect 262 125 263 126
rect 263 125 264 126
rect 265 125 266 126
rect 160 180 161 181
rect 162 180 163 181
rect 163 180 164 181
rect 165 180 166 181
rect 160 181 166 185
rect 160 185 161 186
rect 162 185 163 186
rect 163 185 164 186
rect 165 185 166 186
rect 340 200 341 201
rect 342 200 343 201
rect 343 200 344 201
rect 345 200 346 201
rect 340 201 346 205
rect 340 205 341 206
rect 342 205 343 206
rect 343 205 344 206
rect 345 205 346 206
rect 500 80 501 81
rect 502 80 503 81
rect 503 80 504 81
rect 505 80 506 81
rect 500 81 506 85
rect 500 85 501 86
rect 502 85 503 86
rect 503 85 504 86
rect 505 85 506 86
rect 500 360 501 361
rect 502 360 503 361
rect 503 360 504 361
rect 505 360 506 361
rect 500 361 506 365
rect 500 365 501 366
rect 502 365 503 366
rect 503 365 504 366
rect 505 365 506 366
rect 580 180 581 181
rect 582 180 583 181
rect 583 180 584 181
rect 585 180 586 181
rect 580 181 586 185
rect 580 185 581 186
rect 582 185 583 186
rect 583 185 584 186
rect 585 185 586 186
rect 360 0 361 1
rect 362 0 363 1
rect 363 0 364 1
rect 365 0 366 1
rect 360 1 366 5
rect 360 5 361 6
rect 362 5 363 6
rect 363 5 364 6
rect 365 5 366 6
rect 520 180 521 181
rect 522 180 523 181
rect 523 180 524 181
rect 525 180 526 181
rect 520 181 526 185
rect 520 185 521 186
rect 522 185 523 186
rect 523 185 524 186
rect 525 185 526 186
rect 500 120 501 121
rect 502 120 503 121
rect 503 120 504 121
rect 505 120 506 121
rect 500 121 506 125
rect 500 125 501 126
rect 502 125 503 126
rect 503 125 504 126
rect 505 125 506 126
rect 600 300 601 301
rect 602 300 603 301
rect 603 300 604 301
rect 605 300 606 301
rect 600 301 606 305
rect 600 305 601 306
rect 602 305 603 306
rect 603 305 604 306
rect 605 305 606 306
rect 100 520 101 521
rect 102 520 103 521
rect 103 520 104 521
rect 105 520 106 521
rect 100 521 106 525
rect 100 525 101 526
rect 102 525 103 526
rect 103 525 104 526
rect 105 525 106 526
rect 100 240 101 241
rect 102 240 103 241
rect 103 240 104 241
rect 105 240 106 241
rect 100 241 106 245
rect 100 245 101 246
rect 102 245 103 246
rect 103 245 104 246
rect 105 245 106 246
rect 80 180 81 181
rect 82 180 83 181
rect 83 180 84 181
rect 85 180 86 181
rect 80 181 86 185
rect 80 185 81 186
rect 82 185 83 186
rect 83 185 84 186
rect 85 185 86 186
rect 260 420 261 421
rect 262 420 263 421
rect 263 420 264 421
rect 265 420 266 421
rect 260 421 266 425
rect 260 425 261 426
rect 262 425 263 426
rect 263 425 264 426
rect 265 425 266 426
rect 320 640 321 641
rect 322 640 323 641
rect 323 640 324 641
rect 325 640 326 641
rect 320 641 326 645
rect 320 645 321 646
rect 322 645 323 646
rect 323 645 324 646
rect 325 645 326 646
rect 220 600 221 601
rect 222 600 223 601
rect 223 600 224 601
rect 225 600 226 601
rect 220 601 226 605
rect 220 605 221 606
rect 222 605 223 606
rect 223 605 224 606
rect 225 605 226 606
rect 500 240 501 241
rect 502 240 503 241
rect 503 240 504 241
rect 505 240 506 241
rect 500 241 506 245
rect 500 245 501 246
rect 502 245 503 246
rect 503 245 504 246
rect 505 245 506 246
rect 100 460 101 461
rect 102 460 103 461
rect 103 460 104 461
rect 105 460 106 461
rect 100 461 106 465
rect 100 465 101 466
rect 102 465 103 466
rect 103 465 104 466
rect 105 465 106 466
rect 400 380 401 381
rect 402 380 403 381
rect 403 380 404 381
rect 405 380 406 381
rect 400 381 406 385
rect 400 385 401 386
rect 402 385 403 386
rect 403 385 404 386
rect 405 385 406 386
rect 200 200 201 201
rect 202 200 203 201
rect 203 200 204 201
rect 205 200 206 201
rect 200 201 206 205
rect 200 205 201 206
rect 202 205 203 206
rect 203 205 204 206
rect 205 205 206 206
rect 300 400 301 401
rect 302 400 303 401
rect 303 400 304 401
rect 305 400 306 401
rect 300 401 306 405
rect 300 405 301 406
rect 302 405 303 406
rect 303 405 304 406
rect 305 405 306 406
rect 80 560 81 561
rect 82 560 83 561
rect 83 560 84 561
rect 85 560 86 561
rect 80 561 86 565
rect 80 565 81 566
rect 82 565 83 566
rect 83 565 84 566
rect 85 565 86 566
rect 240 260 241 261
rect 242 260 243 261
rect 243 260 244 261
rect 245 260 246 261
rect 240 261 246 265
rect 240 265 241 266
rect 242 265 243 266
rect 243 265 244 266
rect 245 265 246 266
rect 600 140 601 141
rect 602 140 603 141
rect 603 140 604 141
rect 605 140 606 141
rect 600 141 606 145
rect 600 145 601 146
rect 602 145 603 146
rect 603 145 604 146
rect 605 145 606 146
rect 180 20 181 21
rect 182 20 183 21
rect 183 20 184 21
rect 185 20 186 21
rect 180 21 186 25
rect 180 25 181 26
rect 182 25 183 26
rect 183 25 184 26
rect 185 25 186 26
rect 600 120 601 121
rect 602 120 603 121
rect 603 120 604 121
rect 605 120 606 121
rect 600 121 606 125
rect 600 125 601 126
rect 602 125 603 126
rect 603 125 604 126
rect 605 125 606 126
rect 80 460 81 461
rect 82 460 83 461
rect 83 460 84 461
rect 85 460 86 461
rect 80 461 86 465
rect 80 465 81 466
rect 82 465 83 466
rect 83 465 84 466
rect 85 465 86 466
rect 540 280 541 281
rect 542 280 543 281
rect 543 280 544 281
rect 545 280 546 281
rect 540 281 546 285
rect 540 285 541 286
rect 542 285 543 286
rect 543 285 544 286
rect 545 285 546 286
rect 200 120 201 121
rect 202 120 203 121
rect 203 120 204 121
rect 205 120 206 121
rect 200 121 206 125
rect 200 125 201 126
rect 202 125 203 126
rect 203 125 204 126
rect 205 125 206 126
rect 40 480 41 481
rect 42 480 43 481
rect 43 480 44 481
rect 45 480 46 481
rect 40 481 46 485
rect 40 485 41 486
rect 42 485 43 486
rect 43 485 44 486
rect 45 485 46 486
rect 120 540 121 541
rect 122 540 123 541
rect 123 540 124 541
rect 125 540 126 541
rect 120 541 126 545
rect 120 545 121 546
rect 122 545 123 546
rect 123 545 124 546
rect 125 545 126 546
rect 420 660 421 661
rect 422 660 423 661
rect 423 660 424 661
rect 425 660 426 661
rect 420 661 426 665
rect 420 665 421 666
rect 422 665 423 666
rect 423 665 424 666
rect 425 665 426 666
rect 500 420 501 421
rect 502 420 503 421
rect 503 420 504 421
rect 505 420 506 421
rect 500 421 506 425
rect 500 425 501 426
rect 502 425 503 426
rect 503 425 504 426
rect 505 425 506 426
rect 20 300 21 301
rect 22 300 23 301
rect 23 300 24 301
rect 25 300 26 301
rect 20 301 26 305
rect 20 305 21 306
rect 22 305 23 306
rect 23 305 24 306
rect 25 305 26 306
rect 580 480 581 481
rect 582 480 583 481
rect 583 480 584 481
rect 585 480 586 481
rect 580 481 586 485
rect 580 485 581 486
rect 582 485 583 486
rect 583 485 584 486
rect 585 485 586 486
rect 140 80 141 81
rect 142 80 143 81
rect 143 80 144 81
rect 145 80 146 81
rect 140 81 146 85
rect 140 85 141 86
rect 142 85 143 86
rect 143 85 144 86
rect 145 85 146 86
rect 320 180 321 181
rect 322 180 323 181
rect 323 180 324 181
rect 325 180 326 181
rect 320 181 326 185
rect 320 185 321 186
rect 322 185 323 186
rect 323 185 324 186
rect 325 185 326 186
rect 20 380 21 381
rect 22 380 23 381
rect 23 380 24 381
rect 25 380 26 381
rect 20 381 26 385
rect 20 385 21 386
rect 22 385 23 386
rect 23 385 24 386
rect 25 385 26 386
rect 40 420 41 421
rect 42 420 43 421
rect 43 420 44 421
rect 45 420 46 421
rect 40 421 46 425
rect 40 425 41 426
rect 42 425 43 426
rect 43 425 44 426
rect 45 425 46 426
rect 640 360 641 361
rect 642 360 643 361
rect 643 360 644 361
rect 645 360 646 361
rect 640 361 646 365
rect 640 365 641 366
rect 642 365 643 366
rect 643 365 644 366
rect 645 365 646 366
rect 400 80 401 81
rect 402 80 403 81
rect 403 80 404 81
rect 405 80 406 81
rect 400 81 406 85
rect 400 85 401 86
rect 402 85 403 86
rect 403 85 404 86
rect 405 85 406 86
rect 0 240 1 241
rect 2 240 3 241
rect 3 240 4 241
rect 5 240 6 241
rect 0 241 6 245
rect 0 245 1 246
rect 2 245 3 246
rect 3 245 4 246
rect 5 245 6 246
rect 180 240 181 241
rect 182 240 183 241
rect 183 240 184 241
rect 185 240 186 241
rect 180 241 186 245
rect 180 245 181 246
rect 182 245 183 246
rect 183 245 184 246
rect 185 245 186 246
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect 280 460 281 461
rect 282 460 283 461
rect 283 460 284 461
rect 285 460 286 461
rect 280 461 286 465
rect 280 465 281 466
rect 282 465 283 466
rect 283 465 284 466
rect 285 465 286 466
rect 640 260 641 261
rect 642 260 643 261
rect 643 260 644 261
rect 645 260 646 261
rect 640 261 646 265
rect 640 265 641 266
rect 642 265 643 266
rect 643 265 644 266
rect 645 265 646 266
rect 560 220 561 221
rect 562 220 563 221
rect 563 220 564 221
rect 565 220 566 221
rect 560 221 566 225
rect 560 225 561 226
rect 562 225 563 226
rect 563 225 564 226
rect 565 225 566 226
rect 440 60 441 61
rect 442 60 443 61
rect 443 60 444 61
rect 445 60 446 61
rect 440 61 446 65
rect 440 65 441 66
rect 442 65 443 66
rect 443 65 444 66
rect 445 65 446 66
rect 520 480 521 481
rect 522 480 523 481
rect 523 480 524 481
rect 525 480 526 481
rect 520 481 526 485
rect 520 485 521 486
rect 522 485 523 486
rect 523 485 524 486
rect 525 485 526 486
rect 260 100 261 101
rect 262 100 263 101
rect 263 100 264 101
rect 265 100 266 101
rect 260 101 266 105
rect 260 105 261 106
rect 262 105 263 106
rect 263 105 264 106
rect 265 105 266 106
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect 260 480 261 481
rect 262 480 263 481
rect 263 480 264 481
rect 265 480 266 481
rect 260 481 266 485
rect 260 485 261 486
rect 262 485 263 486
rect 263 485 264 486
rect 265 485 266 486
rect 180 520 181 521
rect 182 520 183 521
rect 183 520 184 521
rect 185 520 186 521
rect 180 521 186 525
rect 180 525 181 526
rect 182 525 183 526
rect 183 525 184 526
rect 185 525 186 526
rect 360 260 361 261
rect 362 260 363 261
rect 363 260 364 261
rect 365 260 366 261
rect 360 261 366 265
rect 360 265 361 266
rect 362 265 363 266
rect 363 265 364 266
rect 365 265 366 266
rect 320 440 321 441
rect 322 440 323 441
rect 323 440 324 441
rect 325 440 326 441
rect 320 441 326 445
rect 320 445 321 446
rect 322 445 323 446
rect 323 445 324 446
rect 325 445 326 446
rect 360 480 361 481
rect 362 480 363 481
rect 363 480 364 481
rect 365 480 366 481
rect 360 481 366 485
rect 360 485 361 486
rect 362 485 363 486
rect 363 485 364 486
rect 365 485 366 486
rect 260 160 261 161
rect 262 160 263 161
rect 263 160 264 161
rect 265 160 266 161
rect 260 161 266 165
rect 260 165 261 166
rect 262 165 263 166
rect 263 165 264 166
rect 265 165 266 166
rect 660 240 661 241
rect 662 240 663 241
rect 663 240 664 241
rect 665 240 666 241
rect 660 241 666 245
rect 660 245 661 246
rect 662 245 663 246
rect 663 245 664 246
rect 665 245 666 246
rect 200 240 201 241
rect 202 240 203 241
rect 203 240 204 241
rect 205 240 206 241
rect 200 241 206 245
rect 200 245 201 246
rect 202 245 203 246
rect 203 245 204 246
rect 205 245 206 246
rect 480 320 481 321
rect 482 320 483 321
rect 483 320 484 321
rect 485 320 486 321
rect 480 321 486 325
rect 480 325 481 326
rect 482 325 483 326
rect 483 325 484 326
rect 485 325 486 326
rect 120 500 121 501
rect 122 500 123 501
rect 123 500 124 501
rect 125 500 126 501
rect 120 501 126 505
rect 120 505 121 506
rect 122 505 123 506
rect 123 505 124 506
rect 125 505 126 506
rect 40 400 41 401
rect 42 400 43 401
rect 43 400 44 401
rect 45 400 46 401
rect 40 401 46 405
rect 40 405 41 406
rect 42 405 43 406
rect 43 405 44 406
rect 45 405 46 406
rect 220 280 221 281
rect 222 280 223 281
rect 223 280 224 281
rect 225 280 226 281
rect 220 281 226 285
rect 220 285 221 286
rect 222 285 223 286
rect 223 285 224 286
rect 225 285 226 286
rect 280 660 281 661
rect 282 660 283 661
rect 283 660 284 661
rect 285 660 286 661
rect 280 661 286 665
rect 280 665 281 666
rect 282 665 283 666
rect 283 665 284 666
rect 285 665 286 666
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect 620 340 621 341
rect 622 340 623 341
rect 623 340 624 341
rect 625 340 626 341
rect 620 341 626 345
rect 620 345 621 346
rect 622 345 623 346
rect 623 345 624 346
rect 625 345 626 346
rect 480 620 481 621
rect 482 620 483 621
rect 483 620 484 621
rect 485 620 486 621
rect 480 621 486 625
rect 480 625 481 626
rect 482 625 483 626
rect 483 625 484 626
rect 485 625 486 626
rect 180 480 181 481
rect 182 480 183 481
rect 183 480 184 481
rect 185 480 186 481
rect 180 481 186 485
rect 180 485 181 486
rect 182 485 183 486
rect 183 485 184 486
rect 185 485 186 486
rect 640 300 641 301
rect 642 300 643 301
rect 643 300 644 301
rect 645 300 646 301
rect 640 301 646 305
rect 640 305 641 306
rect 642 305 643 306
rect 643 305 644 306
rect 645 305 646 306
rect 100 480 101 481
rect 102 480 103 481
rect 103 480 104 481
rect 105 480 106 481
rect 100 481 106 485
rect 100 485 101 486
rect 102 485 103 486
rect 103 485 104 486
rect 105 485 106 486
rect 500 300 501 301
rect 502 300 503 301
rect 503 300 504 301
rect 505 300 506 301
rect 500 301 506 305
rect 500 305 501 306
rect 502 305 503 306
rect 503 305 504 306
rect 505 305 506 306
rect 180 560 181 561
rect 182 560 183 561
rect 183 560 184 561
rect 185 560 186 561
rect 180 561 186 565
rect 180 565 181 566
rect 182 565 183 566
rect 183 565 184 566
rect 185 565 186 566
rect 360 300 361 301
rect 362 300 363 301
rect 363 300 364 301
rect 365 300 366 301
rect 360 301 366 305
rect 360 305 361 306
rect 362 305 363 306
rect 363 305 364 306
rect 365 305 366 306
rect 260 240 261 241
rect 262 240 263 241
rect 263 240 264 241
rect 265 240 266 241
rect 260 241 266 245
rect 260 245 261 246
rect 262 245 263 246
rect 263 245 264 246
rect 265 245 266 246
rect 40 460 41 461
rect 42 460 43 461
rect 43 460 44 461
rect 45 460 46 461
rect 40 461 46 465
rect 40 465 41 466
rect 42 465 43 466
rect 43 465 44 466
rect 45 465 46 466
rect 400 580 401 581
rect 402 580 403 581
rect 403 580 404 581
rect 405 580 406 581
rect 400 581 406 585
rect 400 585 401 586
rect 402 585 403 586
rect 403 585 404 586
rect 405 585 406 586
rect 200 400 201 401
rect 202 400 203 401
rect 203 400 204 401
rect 205 400 206 401
rect 200 401 206 405
rect 200 405 201 406
rect 202 405 203 406
rect 203 405 204 406
rect 205 405 206 406
rect 640 480 641 481
rect 642 480 643 481
rect 643 480 644 481
rect 645 480 646 481
rect 640 481 646 485
rect 640 485 641 486
rect 642 485 643 486
rect 643 485 644 486
rect 645 485 646 486
rect 100 100 101 101
rect 102 100 103 101
rect 103 100 104 101
rect 105 100 106 101
rect 100 101 106 105
rect 100 105 101 106
rect 102 105 103 106
rect 103 105 104 106
rect 105 105 106 106
rect 400 420 401 421
rect 402 420 403 421
rect 403 420 404 421
rect 405 420 406 421
rect 400 421 406 425
rect 400 425 401 426
rect 402 425 403 426
rect 403 425 404 426
rect 405 425 406 426
rect 520 300 521 301
rect 522 300 523 301
rect 523 300 524 301
rect 525 300 526 301
rect 520 301 526 305
rect 520 305 521 306
rect 522 305 523 306
rect 523 305 524 306
rect 525 305 526 306
rect 240 320 241 321
rect 242 320 243 321
rect 243 320 244 321
rect 245 320 246 321
rect 240 321 246 325
rect 240 325 241 326
rect 242 325 243 326
rect 243 325 244 326
rect 245 325 246 326
rect 280 560 281 561
rect 282 560 283 561
rect 283 560 284 561
rect 285 560 286 561
rect 280 561 286 565
rect 280 565 281 566
rect 282 565 283 566
rect 283 565 284 566
rect 285 565 286 566
rect 40 440 41 441
rect 42 440 43 441
rect 43 440 44 441
rect 45 440 46 441
rect 40 441 46 445
rect 40 445 41 446
rect 42 445 43 446
rect 43 445 44 446
rect 45 445 46 446
rect 0 160 1 161
rect 2 160 3 161
rect 3 160 4 161
rect 5 160 6 161
rect 0 161 6 165
rect 0 165 1 166
rect 2 165 3 166
rect 3 165 4 166
rect 5 165 6 166
rect 260 180 261 181
rect 262 180 263 181
rect 263 180 264 181
rect 265 180 266 181
rect 260 181 266 185
rect 260 185 261 186
rect 262 185 263 186
rect 263 185 264 186
rect 265 185 266 186
rect 400 460 401 461
rect 402 460 403 461
rect 403 460 404 461
rect 405 460 406 461
rect 400 461 406 465
rect 400 465 401 466
rect 402 465 403 466
rect 403 465 404 466
rect 405 465 406 466
rect 600 380 601 381
rect 602 380 603 381
rect 603 380 604 381
rect 605 380 606 381
rect 600 381 606 385
rect 600 385 601 386
rect 602 385 603 386
rect 603 385 604 386
rect 605 385 606 386
rect 160 220 161 221
rect 162 220 163 221
rect 163 220 164 221
rect 165 220 166 221
rect 160 221 166 225
rect 160 225 161 226
rect 162 225 163 226
rect 163 225 164 226
rect 165 225 166 226
rect 220 560 221 561
rect 222 560 223 561
rect 223 560 224 561
rect 225 560 226 561
rect 220 561 226 565
rect 220 565 221 566
rect 222 565 223 566
rect 223 565 224 566
rect 225 565 226 566
rect 480 160 481 161
rect 482 160 483 161
rect 483 160 484 161
rect 485 160 486 161
rect 480 161 486 165
rect 480 165 481 166
rect 482 165 483 166
rect 483 165 484 166
rect 485 165 486 166
rect 300 500 301 501
rect 302 500 303 501
rect 303 500 304 501
rect 305 500 306 501
rect 300 501 306 505
rect 300 505 301 506
rect 302 505 303 506
rect 303 505 304 506
rect 305 505 306 506
rect 80 400 81 401
rect 82 400 83 401
rect 83 400 84 401
rect 85 400 86 401
rect 80 401 86 405
rect 80 405 81 406
rect 82 405 83 406
rect 83 405 84 406
rect 85 405 86 406
rect 340 340 341 341
rect 342 340 343 341
rect 343 340 344 341
rect 345 340 346 341
rect 340 341 346 345
rect 340 345 341 346
rect 342 345 343 346
rect 343 345 344 346
rect 345 345 346 346
rect 400 0 401 1
rect 402 0 403 1
rect 403 0 404 1
rect 405 0 406 1
rect 400 1 406 5
rect 400 5 401 6
rect 402 5 403 6
rect 403 5 404 6
rect 405 5 406 6
rect 480 180 481 181
rect 482 180 483 181
rect 483 180 484 181
rect 485 180 486 181
rect 480 181 486 185
rect 480 185 481 186
rect 482 185 483 186
rect 483 185 484 186
rect 485 185 486 186
rect 420 400 421 401
rect 422 400 423 401
rect 423 400 424 401
rect 425 400 426 401
rect 420 401 426 405
rect 420 405 421 406
rect 422 405 423 406
rect 423 405 424 406
rect 425 405 426 406
rect 280 580 281 581
rect 282 580 283 581
rect 283 580 284 581
rect 285 580 286 581
rect 280 581 286 585
rect 280 585 281 586
rect 282 585 283 586
rect 283 585 284 586
rect 285 585 286 586
rect 440 120 441 121
rect 442 120 443 121
rect 443 120 444 121
rect 445 120 446 121
rect 440 121 446 125
rect 440 125 441 126
rect 442 125 443 126
rect 443 125 444 126
rect 445 125 446 126
rect 180 60 181 61
rect 182 60 183 61
rect 183 60 184 61
rect 185 60 186 61
rect 180 61 186 65
rect 180 65 181 66
rect 182 65 183 66
rect 183 65 184 66
rect 185 65 186 66
rect 460 400 461 401
rect 462 400 463 401
rect 463 400 464 401
rect 465 400 466 401
rect 460 401 466 405
rect 460 405 461 406
rect 462 405 463 406
rect 463 405 464 406
rect 465 405 466 406
rect 560 400 561 401
rect 562 400 563 401
rect 563 400 564 401
rect 565 400 566 401
rect 560 401 566 405
rect 560 405 561 406
rect 562 405 563 406
rect 563 405 564 406
rect 565 405 566 406
rect 540 140 541 141
rect 542 140 543 141
rect 543 140 544 141
rect 545 140 546 141
rect 540 141 546 145
rect 540 145 541 146
rect 542 145 543 146
rect 543 145 544 146
rect 545 145 546 146
rect 180 380 181 381
rect 182 380 183 381
rect 183 380 184 381
rect 185 380 186 381
rect 180 381 186 385
rect 180 385 181 386
rect 182 385 183 386
rect 183 385 184 386
rect 185 385 186 386
rect 600 440 601 441
rect 602 440 603 441
rect 603 440 604 441
rect 605 440 606 441
rect 600 441 606 445
rect 600 445 601 446
rect 602 445 603 446
rect 603 445 604 446
rect 605 445 606 446
rect 480 100 481 101
rect 482 100 483 101
rect 483 100 484 101
rect 485 100 486 101
rect 480 101 486 105
rect 480 105 481 106
rect 482 105 483 106
rect 483 105 484 106
rect 485 105 486 106
rect 240 520 241 521
rect 242 520 243 521
rect 243 520 244 521
rect 245 520 246 521
rect 240 521 246 525
rect 240 525 241 526
rect 242 525 243 526
rect 243 525 244 526
rect 245 525 246 526
rect 240 580 241 581
rect 242 580 243 581
rect 243 580 244 581
rect 245 580 246 581
rect 240 581 246 585
rect 240 585 241 586
rect 242 585 243 586
rect 243 585 244 586
rect 245 585 246 586
rect 380 180 381 181
rect 382 180 383 181
rect 383 180 384 181
rect 385 180 386 181
rect 380 181 386 185
rect 380 185 381 186
rect 382 185 383 186
rect 383 185 384 186
rect 385 185 386 186
rect 640 380 641 381
rect 642 380 643 381
rect 643 380 644 381
rect 645 380 646 381
rect 640 381 646 385
rect 640 385 641 386
rect 642 385 643 386
rect 643 385 644 386
rect 645 385 646 386
rect 340 500 341 501
rect 342 500 343 501
rect 343 500 344 501
rect 345 500 346 501
rect 340 501 346 505
rect 340 505 341 506
rect 342 505 343 506
rect 343 505 344 506
rect 345 505 346 506
rect 60 500 61 501
rect 62 500 63 501
rect 63 500 64 501
rect 65 500 66 501
rect 60 501 66 505
rect 60 505 61 506
rect 62 505 63 506
rect 63 505 64 506
rect 65 505 66 506
rect 200 320 201 321
rect 202 320 203 321
rect 203 320 204 321
rect 205 320 206 321
rect 200 321 206 325
rect 200 325 201 326
rect 202 325 203 326
rect 203 325 204 326
rect 205 325 206 326
rect 580 160 581 161
rect 582 160 583 161
rect 583 160 584 161
rect 585 160 586 161
rect 580 161 586 165
rect 580 165 581 166
rect 582 165 583 166
rect 583 165 584 166
rect 585 165 586 166
rect 120 80 121 81
rect 122 80 123 81
rect 123 80 124 81
rect 125 80 126 81
rect 120 81 126 85
rect 120 85 121 86
rect 122 85 123 86
rect 123 85 124 86
rect 125 85 126 86
rect 440 540 441 541
rect 442 540 443 541
rect 443 540 444 541
rect 445 540 446 541
rect 440 541 446 545
rect 440 545 441 546
rect 442 545 443 546
rect 443 545 444 546
rect 445 545 446 546
rect 140 60 141 61
rect 142 60 143 61
rect 143 60 144 61
rect 145 60 146 61
rect 140 61 146 65
rect 140 65 141 66
rect 142 65 143 66
rect 143 65 144 66
rect 145 65 146 66
rect 0 460 1 461
rect 2 460 3 461
rect 3 460 4 461
rect 5 460 6 461
rect 0 461 6 465
rect 0 465 1 466
rect 2 465 3 466
rect 3 465 4 466
rect 5 465 6 466
rect 620 280 621 281
rect 622 280 623 281
rect 623 280 624 281
rect 625 280 626 281
rect 620 281 626 285
rect 620 285 621 286
rect 622 285 623 286
rect 623 285 624 286
rect 625 285 626 286
rect 480 560 481 561
rect 482 560 483 561
rect 483 560 484 561
rect 485 560 486 561
rect 480 561 486 565
rect 480 565 481 566
rect 482 565 483 566
rect 483 565 484 566
rect 485 565 486 566
rect 20 460 21 461
rect 22 460 23 461
rect 23 460 24 461
rect 25 460 26 461
rect 20 461 26 465
rect 20 465 21 466
rect 22 465 23 466
rect 23 465 24 466
rect 25 465 26 466
rect 480 260 481 261
rect 482 260 483 261
rect 483 260 484 261
rect 485 260 486 261
rect 480 261 486 265
rect 480 265 481 266
rect 482 265 483 266
rect 483 265 484 266
rect 485 265 486 266
rect 260 540 261 541
rect 262 540 263 541
rect 263 540 264 541
rect 265 540 266 541
rect 260 541 266 545
rect 260 545 261 546
rect 262 545 263 546
rect 263 545 264 546
rect 265 545 266 546
rect 260 0 261 1
rect 262 0 263 1
rect 263 0 264 1
rect 265 0 266 1
rect 260 1 266 5
rect 260 5 261 6
rect 262 5 263 6
rect 263 5 264 6
rect 265 5 266 6
rect 80 260 81 261
rect 82 260 83 261
rect 83 260 84 261
rect 85 260 86 261
rect 80 261 86 265
rect 80 265 81 266
rect 82 265 83 266
rect 83 265 84 266
rect 85 265 86 266
rect 480 480 481 481
rect 482 480 483 481
rect 483 480 484 481
rect 485 480 486 481
rect 480 481 486 485
rect 480 485 481 486
rect 482 485 483 486
rect 483 485 484 486
rect 485 485 486 486
rect 280 240 281 241
rect 282 240 283 241
rect 283 240 284 241
rect 285 240 286 241
rect 280 241 286 245
rect 280 245 281 246
rect 282 245 283 246
rect 283 245 284 246
rect 285 245 286 246
rect 460 640 461 641
rect 462 640 463 641
rect 463 640 464 641
rect 465 640 466 641
rect 460 641 466 645
rect 460 645 461 646
rect 462 645 463 646
rect 463 645 464 646
rect 465 645 466 646
rect 460 460 461 461
rect 462 460 463 461
rect 463 460 464 461
rect 465 460 466 461
rect 460 461 466 465
rect 460 465 461 466
rect 462 465 463 466
rect 463 465 464 466
rect 465 465 466 466
rect 340 360 341 361
rect 342 360 343 361
rect 343 360 344 361
rect 345 360 346 361
rect 340 361 346 365
rect 340 365 341 366
rect 342 365 343 366
rect 343 365 344 366
rect 345 365 346 366
rect 300 140 301 141
rect 302 140 303 141
rect 303 140 304 141
rect 305 140 306 141
rect 300 141 306 145
rect 300 145 301 146
rect 302 145 303 146
rect 303 145 304 146
rect 305 145 306 146
rect 660 260 661 261
rect 662 260 663 261
rect 663 260 664 261
rect 665 260 666 261
rect 660 261 666 265
rect 660 265 661 266
rect 662 265 663 266
rect 663 265 664 266
rect 665 265 666 266
rect 380 260 381 261
rect 382 260 383 261
rect 383 260 384 261
rect 385 260 386 261
rect 380 261 386 265
rect 380 265 381 266
rect 382 265 383 266
rect 383 265 384 266
rect 385 265 386 266
rect 80 60 81 61
rect 82 60 83 61
rect 83 60 84 61
rect 85 60 86 61
rect 80 61 86 65
rect 80 65 81 66
rect 82 65 83 66
rect 83 65 84 66
rect 85 65 86 66
rect 340 300 341 301
rect 342 300 343 301
rect 343 300 344 301
rect 345 300 346 301
rect 340 301 346 305
rect 340 305 341 306
rect 342 305 343 306
rect 343 305 344 306
rect 345 305 346 306
rect 160 600 161 601
rect 162 600 163 601
rect 163 600 164 601
rect 165 600 166 601
rect 160 601 166 605
rect 160 605 161 606
rect 162 605 163 606
rect 163 605 164 606
rect 165 605 166 606
rect 340 20 341 21
rect 342 20 343 21
rect 343 20 344 21
rect 345 20 346 21
rect 340 21 346 25
rect 340 25 341 26
rect 342 25 343 26
rect 343 25 344 26
rect 345 25 346 26
rect 300 460 301 461
rect 302 460 303 461
rect 303 460 304 461
rect 305 460 306 461
rect 300 461 306 465
rect 300 465 301 466
rect 302 465 303 466
rect 303 465 304 466
rect 305 465 306 466
rect 180 0 181 1
rect 182 0 183 1
rect 183 0 184 1
rect 185 0 186 1
rect 180 1 186 5
rect 180 5 181 6
rect 182 5 183 6
rect 183 5 184 6
rect 185 5 186 6
rect 100 560 101 561
rect 102 560 103 561
rect 103 560 104 561
rect 105 560 106 561
rect 100 561 106 565
rect 100 565 101 566
rect 102 565 103 566
rect 103 565 104 566
rect 105 565 106 566
rect 380 80 381 81
rect 382 80 383 81
rect 383 80 384 81
rect 385 80 386 81
rect 380 81 386 85
rect 380 85 381 86
rect 382 85 383 86
rect 383 85 384 86
rect 385 85 386 86
rect 420 0 421 1
rect 422 0 423 1
rect 423 0 424 1
rect 425 0 426 1
rect 420 1 426 5
rect 420 5 421 6
rect 422 5 423 6
rect 423 5 424 6
rect 425 5 426 6
rect 560 440 561 441
rect 562 440 563 441
rect 563 440 564 441
rect 565 440 566 441
rect 560 441 566 445
rect 560 445 561 446
rect 562 445 563 446
rect 563 445 564 446
rect 565 445 566 446
rect 440 480 441 481
rect 442 480 443 481
rect 443 480 444 481
rect 445 480 446 481
rect 440 481 446 485
rect 440 485 441 486
rect 442 485 443 486
rect 443 485 444 486
rect 445 485 446 486
rect 300 20 301 21
rect 302 20 303 21
rect 303 20 304 21
rect 305 20 306 21
rect 300 21 306 25
rect 300 25 301 26
rect 302 25 303 26
rect 303 25 304 26
rect 305 25 306 26
rect 20 140 21 141
rect 22 140 23 141
rect 23 140 24 141
rect 25 140 26 141
rect 20 141 26 145
rect 20 145 21 146
rect 22 145 23 146
rect 23 145 24 146
rect 25 145 26 146
rect 100 40 101 41
rect 102 40 103 41
rect 103 40 104 41
rect 105 40 106 41
rect 100 41 106 45
rect 100 45 101 46
rect 102 45 103 46
rect 103 45 104 46
rect 105 45 106 46
rect 520 160 521 161
rect 522 160 523 161
rect 523 160 524 161
rect 525 160 526 161
rect 520 161 526 165
rect 520 165 521 166
rect 522 165 523 166
rect 523 165 524 166
rect 525 165 526 166
rect 340 620 341 621
rect 342 620 343 621
rect 343 620 344 621
rect 345 620 346 621
rect 340 621 346 625
rect 340 625 341 626
rect 342 625 343 626
rect 343 625 344 626
rect 345 625 346 626
rect 540 260 541 261
rect 542 260 543 261
rect 543 260 544 261
rect 545 260 546 261
rect 540 261 546 265
rect 540 265 541 266
rect 542 265 543 266
rect 543 265 544 266
rect 545 265 546 266
rect 420 260 421 261
rect 422 260 423 261
rect 423 260 424 261
rect 425 260 426 261
rect 420 261 426 265
rect 420 265 421 266
rect 422 265 423 266
rect 423 265 424 266
rect 425 265 426 266
rect 640 460 641 461
rect 642 460 643 461
rect 643 460 644 461
rect 645 460 646 461
rect 640 461 646 465
rect 640 465 641 466
rect 642 465 643 466
rect 643 465 644 466
rect 645 465 646 466
rect 460 320 461 321
rect 462 320 463 321
rect 463 320 464 321
rect 465 320 466 321
rect 460 321 466 325
rect 460 325 461 326
rect 462 325 463 326
rect 463 325 464 326
rect 465 325 466 326
rect 300 0 301 1
rect 302 0 303 1
rect 303 0 304 1
rect 305 0 306 1
rect 300 1 306 5
rect 300 5 301 6
rect 302 5 303 6
rect 303 5 304 6
rect 305 5 306 6
rect 60 320 61 321
rect 62 320 63 321
rect 63 320 64 321
rect 65 320 66 321
rect 60 321 66 325
rect 60 325 61 326
rect 62 325 63 326
rect 63 325 64 326
rect 65 325 66 326
rect 300 560 301 561
rect 302 560 303 561
rect 303 560 304 561
rect 305 560 306 561
rect 300 561 306 565
rect 300 565 301 566
rect 302 565 303 566
rect 303 565 304 566
rect 305 565 306 566
rect 80 320 81 321
rect 82 320 83 321
rect 83 320 84 321
rect 85 320 86 321
rect 80 321 86 325
rect 80 325 81 326
rect 82 325 83 326
rect 83 325 84 326
rect 85 325 86 326
rect 100 200 101 201
rect 102 200 103 201
rect 103 200 104 201
rect 105 200 106 201
rect 100 201 106 205
rect 100 205 101 206
rect 102 205 103 206
rect 103 205 104 206
rect 105 205 106 206
rect 160 320 161 321
rect 162 320 163 321
rect 163 320 164 321
rect 165 320 166 321
rect 160 321 166 325
rect 160 325 161 326
rect 162 325 163 326
rect 163 325 164 326
rect 165 325 166 326
rect 400 300 401 301
rect 402 300 403 301
rect 403 300 404 301
rect 405 300 406 301
rect 400 301 406 305
rect 400 305 401 306
rect 402 305 403 306
rect 403 305 404 306
rect 405 305 406 306
rect 400 480 401 481
rect 402 480 403 481
rect 403 480 404 481
rect 405 480 406 481
rect 400 481 406 485
rect 400 485 401 486
rect 402 485 403 486
rect 403 485 404 486
rect 405 485 406 486
rect 60 380 61 381
rect 62 380 63 381
rect 63 380 64 381
rect 65 380 66 381
rect 60 381 66 385
rect 60 385 61 386
rect 62 385 63 386
rect 63 385 64 386
rect 65 385 66 386
rect 140 540 141 541
rect 142 540 143 541
rect 143 540 144 541
rect 145 540 146 541
rect 140 541 146 545
rect 140 545 141 546
rect 142 545 143 546
rect 143 545 144 546
rect 145 545 146 546
rect 200 600 201 601
rect 202 600 203 601
rect 203 600 204 601
rect 205 600 206 601
rect 200 601 206 605
rect 200 605 201 606
rect 202 605 203 606
rect 203 605 204 606
rect 205 605 206 606
rect 220 480 221 481
rect 222 480 223 481
rect 223 480 224 481
rect 225 480 226 481
rect 220 481 226 485
rect 220 485 221 486
rect 222 485 223 486
rect 223 485 224 486
rect 225 485 226 486
rect 140 240 141 241
rect 142 240 143 241
rect 143 240 144 241
rect 145 240 146 241
rect 140 241 146 245
rect 140 245 141 246
rect 142 245 143 246
rect 143 245 144 246
rect 145 245 146 246
rect 140 20 141 21
rect 142 20 143 21
rect 143 20 144 21
rect 145 20 146 21
rect 140 21 146 25
rect 140 25 141 26
rect 142 25 143 26
rect 143 25 144 26
rect 145 25 146 26
rect 200 60 201 61
rect 202 60 203 61
rect 203 60 204 61
rect 205 60 206 61
rect 200 61 206 65
rect 200 65 201 66
rect 202 65 203 66
rect 203 65 204 66
rect 205 65 206 66
rect 240 280 241 281
rect 242 280 243 281
rect 243 280 244 281
rect 245 280 246 281
rect 240 281 246 285
rect 240 285 241 286
rect 242 285 243 286
rect 243 285 244 286
rect 245 285 246 286
rect 360 240 361 241
rect 362 240 363 241
rect 363 240 364 241
rect 365 240 366 241
rect 360 241 366 245
rect 360 245 361 246
rect 362 245 363 246
rect 363 245 364 246
rect 365 245 366 246
rect 480 140 481 141
rect 482 140 483 141
rect 483 140 484 141
rect 485 140 486 141
rect 480 141 486 145
rect 480 145 481 146
rect 482 145 483 146
rect 483 145 484 146
rect 485 145 486 146
rect 220 580 221 581
rect 222 580 223 581
rect 223 580 224 581
rect 225 580 226 581
rect 220 581 226 585
rect 220 585 221 586
rect 222 585 223 586
rect 223 585 224 586
rect 225 585 226 586
rect 220 460 221 461
rect 222 460 223 461
rect 223 460 224 461
rect 225 460 226 461
rect 220 461 226 465
rect 220 465 221 466
rect 222 465 223 466
rect 223 465 224 466
rect 225 465 226 466
rect 240 420 241 421
rect 242 420 243 421
rect 243 420 244 421
rect 245 420 246 421
rect 240 421 246 425
rect 240 425 241 426
rect 242 425 243 426
rect 243 425 244 426
rect 245 425 246 426
rect 180 220 181 221
rect 182 220 183 221
rect 183 220 184 221
rect 185 220 186 221
rect 180 221 186 225
rect 180 225 181 226
rect 182 225 183 226
rect 183 225 184 226
rect 185 225 186 226
rect 380 620 381 621
rect 382 620 383 621
rect 383 620 384 621
rect 385 620 386 621
rect 380 621 386 625
rect 380 625 381 626
rect 382 625 383 626
rect 383 625 384 626
rect 385 625 386 626
rect 0 220 1 221
rect 2 220 3 221
rect 3 220 4 221
rect 5 220 6 221
rect 0 221 6 225
rect 0 225 1 226
rect 2 225 3 226
rect 3 225 4 226
rect 5 225 6 226
rect 560 460 561 461
rect 562 460 563 461
rect 563 460 564 461
rect 565 460 566 461
rect 560 461 566 465
rect 560 465 561 466
rect 562 465 563 466
rect 563 465 564 466
rect 565 465 566 466
rect 320 340 321 341
rect 322 340 323 341
rect 323 340 324 341
rect 325 340 326 341
rect 320 341 326 345
rect 320 345 321 346
rect 322 345 323 346
rect 323 345 324 346
rect 325 345 326 346
rect 40 300 41 301
rect 42 300 43 301
rect 43 300 44 301
rect 45 300 46 301
rect 40 301 46 305
rect 40 305 41 306
rect 42 305 43 306
rect 43 305 44 306
rect 45 305 46 306
rect 600 340 601 341
rect 602 340 603 341
rect 603 340 604 341
rect 605 340 606 341
rect 600 341 606 345
rect 600 345 601 346
rect 602 345 603 346
rect 603 345 604 346
rect 605 345 606 346
rect 280 600 281 601
rect 282 600 283 601
rect 283 600 284 601
rect 285 600 286 601
rect 280 601 286 605
rect 280 605 281 606
rect 282 605 283 606
rect 283 605 284 606
rect 285 605 286 606
rect 580 320 581 321
rect 582 320 583 321
rect 583 320 584 321
rect 585 320 586 321
rect 580 321 586 325
rect 580 325 581 326
rect 582 325 583 326
rect 583 325 584 326
rect 585 325 586 326
rect 460 0 461 1
rect 462 0 463 1
rect 463 0 464 1
rect 465 0 466 1
rect 460 1 466 5
rect 460 5 461 6
rect 462 5 463 6
rect 463 5 464 6
rect 465 5 466 6
rect 240 500 241 501
rect 242 500 243 501
rect 243 500 244 501
rect 245 500 246 501
rect 240 501 246 505
rect 240 505 241 506
rect 242 505 243 506
rect 243 505 244 506
rect 245 505 246 506
rect 320 620 321 621
rect 322 620 323 621
rect 323 620 324 621
rect 325 620 326 621
rect 320 621 326 625
rect 320 625 321 626
rect 322 625 323 626
rect 323 625 324 626
rect 325 625 326 626
rect 480 520 481 521
rect 482 520 483 521
rect 483 520 484 521
rect 485 520 486 521
rect 480 521 486 525
rect 480 525 481 526
rect 482 525 483 526
rect 483 525 484 526
rect 485 525 486 526
rect 400 280 401 281
rect 402 280 403 281
rect 403 280 404 281
rect 405 280 406 281
rect 400 281 406 285
rect 400 285 401 286
rect 402 285 403 286
rect 403 285 404 286
rect 405 285 406 286
rect 420 560 421 561
rect 422 560 423 561
rect 423 560 424 561
rect 425 560 426 561
rect 420 561 426 565
rect 420 565 421 566
rect 422 565 423 566
rect 423 565 424 566
rect 425 565 426 566
rect 160 400 161 401
rect 162 400 163 401
rect 163 400 164 401
rect 165 400 166 401
rect 160 401 166 405
rect 160 405 161 406
rect 162 405 163 406
rect 163 405 164 406
rect 165 405 166 406
rect 400 60 401 61
rect 402 60 403 61
rect 403 60 404 61
rect 405 60 406 61
rect 400 61 406 65
rect 400 65 401 66
rect 402 65 403 66
rect 403 65 404 66
rect 405 65 406 66
rect 580 100 581 101
rect 582 100 583 101
rect 583 100 584 101
rect 585 100 586 101
rect 580 101 586 105
rect 580 105 581 106
rect 582 105 583 106
rect 583 105 584 106
rect 585 105 586 106
rect 180 300 181 301
rect 182 300 183 301
rect 183 300 184 301
rect 185 300 186 301
rect 180 301 186 305
rect 180 305 181 306
rect 182 305 183 306
rect 183 305 184 306
rect 185 305 186 306
rect 0 320 1 321
rect 2 320 3 321
rect 3 320 4 321
rect 5 320 6 321
rect 0 321 6 325
rect 0 325 1 326
rect 2 325 3 326
rect 3 325 4 326
rect 5 325 6 326
rect 120 240 121 241
rect 122 240 123 241
rect 123 240 124 241
rect 125 240 126 241
rect 120 241 126 245
rect 120 245 121 246
rect 122 245 123 246
rect 123 245 124 246
rect 125 245 126 246
rect 420 20 421 21
rect 422 20 423 21
rect 423 20 424 21
rect 425 20 426 21
rect 420 21 426 25
rect 420 25 421 26
rect 422 25 423 26
rect 423 25 424 26
rect 425 25 426 26
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect 160 20 161 21
rect 162 20 163 21
rect 163 20 164 21
rect 165 20 166 21
rect 160 21 166 25
rect 160 25 161 26
rect 162 25 163 26
rect 163 25 164 26
rect 165 25 166 26
rect 520 520 521 521
rect 522 520 523 521
rect 523 520 524 521
rect 525 520 526 521
rect 520 521 526 525
rect 520 525 521 526
rect 522 525 523 526
rect 523 525 524 526
rect 525 525 526 526
rect 260 600 261 601
rect 262 600 263 601
rect 263 600 264 601
rect 265 600 266 601
rect 260 601 266 605
rect 260 605 261 606
rect 262 605 263 606
rect 263 605 264 606
rect 265 605 266 606
rect 560 540 561 541
rect 562 540 563 541
rect 563 540 564 541
rect 565 540 566 541
rect 560 541 566 545
rect 560 545 561 546
rect 562 545 563 546
rect 563 545 564 546
rect 565 545 566 546
rect 140 400 141 401
rect 142 400 143 401
rect 143 400 144 401
rect 145 400 146 401
rect 140 401 146 405
rect 140 405 141 406
rect 142 405 143 406
rect 143 405 144 406
rect 145 405 146 406
rect 400 620 401 621
rect 402 620 403 621
rect 403 620 404 621
rect 405 620 406 621
rect 400 621 406 625
rect 400 625 401 626
rect 402 625 403 626
rect 403 625 404 626
rect 405 625 406 626
rect 640 240 641 241
rect 642 240 643 241
rect 643 240 644 241
rect 645 240 646 241
rect 640 241 646 245
rect 640 245 641 246
rect 642 245 643 246
rect 643 245 644 246
rect 645 245 646 246
rect 540 240 541 241
rect 542 240 543 241
rect 543 240 544 241
rect 545 240 546 241
rect 540 241 546 245
rect 540 245 541 246
rect 542 245 543 246
rect 543 245 544 246
rect 545 245 546 246
rect 460 480 461 481
rect 462 480 463 481
rect 463 480 464 481
rect 465 480 466 481
rect 460 481 466 485
rect 460 485 461 486
rect 462 485 463 486
rect 463 485 464 486
rect 465 485 466 486
rect 20 520 21 521
rect 22 520 23 521
rect 23 520 24 521
rect 25 520 26 521
rect 20 521 26 525
rect 20 525 21 526
rect 22 525 23 526
rect 23 525 24 526
rect 25 525 26 526
rect 440 40 441 41
rect 442 40 443 41
rect 443 40 444 41
rect 445 40 446 41
rect 440 41 446 45
rect 440 45 441 46
rect 442 45 443 46
rect 443 45 444 46
rect 445 45 446 46
rect 460 360 461 361
rect 462 360 463 361
rect 463 360 464 361
rect 465 360 466 361
rect 460 361 466 365
rect 460 365 461 366
rect 462 365 463 366
rect 463 365 464 366
rect 465 365 466 366
rect 60 520 61 521
rect 62 520 63 521
rect 63 520 64 521
rect 65 520 66 521
rect 60 521 66 525
rect 60 525 61 526
rect 62 525 63 526
rect 63 525 64 526
rect 65 525 66 526
rect 340 440 341 441
rect 342 440 343 441
rect 343 440 344 441
rect 345 440 346 441
rect 340 441 346 445
rect 340 445 341 446
rect 342 445 343 446
rect 343 445 344 446
rect 345 445 346 446
rect 380 120 381 121
rect 382 120 383 121
rect 383 120 384 121
rect 385 120 386 121
rect 380 121 386 125
rect 380 125 381 126
rect 382 125 383 126
rect 383 125 384 126
rect 385 125 386 126
rect 80 580 81 581
rect 82 580 83 581
rect 83 580 84 581
rect 85 580 86 581
rect 80 581 86 585
rect 80 585 81 586
rect 82 585 83 586
rect 83 585 84 586
rect 85 585 86 586
rect 580 340 581 341
rect 582 340 583 341
rect 583 340 584 341
rect 585 340 586 341
rect 580 341 586 345
rect 580 345 581 346
rect 582 345 583 346
rect 583 345 584 346
rect 585 345 586 346
rect 360 220 361 221
rect 362 220 363 221
rect 363 220 364 221
rect 365 220 366 221
rect 360 221 366 225
rect 360 225 361 226
rect 362 225 363 226
rect 363 225 364 226
rect 365 225 366 226
rect 440 100 441 101
rect 442 100 443 101
rect 443 100 444 101
rect 445 100 446 101
rect 440 101 446 105
rect 440 105 441 106
rect 442 105 443 106
rect 443 105 444 106
rect 445 105 446 106
rect 80 340 81 341
rect 82 340 83 341
rect 83 340 84 341
rect 85 340 86 341
rect 80 341 86 345
rect 80 345 81 346
rect 82 345 83 346
rect 83 345 84 346
rect 85 345 86 346
rect 120 20 121 21
rect 122 20 123 21
rect 123 20 124 21
rect 125 20 126 21
rect 120 21 126 25
rect 120 25 121 26
rect 122 25 123 26
rect 123 25 124 26
rect 125 25 126 26
rect 300 600 301 601
rect 302 600 303 601
rect 303 600 304 601
rect 305 600 306 601
rect 300 601 306 605
rect 300 605 301 606
rect 302 605 303 606
rect 303 605 304 606
rect 305 605 306 606
rect 180 100 181 101
rect 182 100 183 101
rect 183 100 184 101
rect 185 100 186 101
rect 180 101 186 105
rect 180 105 181 106
rect 182 105 183 106
rect 183 105 184 106
rect 185 105 186 106
rect 660 200 661 201
rect 662 200 663 201
rect 663 200 664 201
rect 665 200 666 201
rect 660 201 666 205
rect 660 205 661 206
rect 662 205 663 206
rect 663 205 664 206
rect 665 205 666 206
rect 20 260 21 261
rect 22 260 23 261
rect 23 260 24 261
rect 25 260 26 261
rect 20 261 26 265
rect 20 265 21 266
rect 22 265 23 266
rect 23 265 24 266
rect 25 265 26 266
rect 380 300 381 301
rect 382 300 383 301
rect 383 300 384 301
rect 385 300 386 301
rect 380 301 386 305
rect 380 305 381 306
rect 382 305 383 306
rect 383 305 384 306
rect 385 305 386 306
rect 400 240 401 241
rect 402 240 403 241
rect 403 240 404 241
rect 405 240 406 241
rect 400 241 406 245
rect 400 245 401 246
rect 402 245 403 246
rect 403 245 404 246
rect 405 245 406 246
rect 60 300 61 301
rect 62 300 63 301
rect 63 300 64 301
rect 65 300 66 301
rect 60 301 66 305
rect 60 305 61 306
rect 62 305 63 306
rect 63 305 64 306
rect 65 305 66 306
rect 580 520 581 521
rect 582 520 583 521
rect 583 520 584 521
rect 585 520 586 521
rect 580 521 586 525
rect 580 525 581 526
rect 582 525 583 526
rect 583 525 584 526
rect 585 525 586 526
rect 420 620 421 621
rect 422 620 423 621
rect 423 620 424 621
rect 425 620 426 621
rect 420 621 426 625
rect 420 625 421 626
rect 422 625 423 626
rect 423 625 424 626
rect 425 625 426 626
rect 20 200 21 201
rect 22 200 23 201
rect 23 200 24 201
rect 25 200 26 201
rect 20 201 26 205
rect 20 205 21 206
rect 22 205 23 206
rect 23 205 24 206
rect 25 205 26 206
rect 500 260 501 261
rect 502 260 503 261
rect 503 260 504 261
rect 505 260 506 261
rect 500 261 506 265
rect 500 265 501 266
rect 502 265 503 266
rect 503 265 504 266
rect 505 265 506 266
rect 260 220 261 221
rect 262 220 263 221
rect 263 220 264 221
rect 265 220 266 221
rect 260 221 266 225
rect 260 225 261 226
rect 262 225 263 226
rect 263 225 264 226
rect 265 225 266 226
rect 80 280 81 281
rect 82 280 83 281
rect 83 280 84 281
rect 85 280 86 281
rect 80 281 86 285
rect 80 285 81 286
rect 82 285 83 286
rect 83 285 84 286
rect 85 285 86 286
rect 160 140 161 141
rect 162 140 163 141
rect 163 140 164 141
rect 165 140 166 141
rect 160 141 166 145
rect 160 145 161 146
rect 162 145 163 146
rect 163 145 164 146
rect 165 145 166 146
rect 220 420 221 421
rect 222 420 223 421
rect 223 420 224 421
rect 225 420 226 421
rect 220 421 226 425
rect 220 425 221 426
rect 222 425 223 426
rect 223 425 224 426
rect 225 425 226 426
rect 120 200 121 201
rect 122 200 123 201
rect 123 200 124 201
rect 125 200 126 201
rect 120 201 126 205
rect 120 205 121 206
rect 122 205 123 206
rect 123 205 124 206
rect 125 205 126 206
rect 360 620 361 621
rect 362 620 363 621
rect 363 620 364 621
rect 365 620 366 621
rect 360 621 366 625
rect 360 625 361 626
rect 362 625 363 626
rect 363 625 364 626
rect 365 625 366 626
rect 620 260 621 261
rect 622 260 623 261
rect 623 260 624 261
rect 625 260 626 261
rect 620 261 626 265
rect 620 265 621 266
rect 622 265 623 266
rect 623 265 624 266
rect 625 265 626 266
rect 60 200 61 201
rect 62 200 63 201
rect 63 200 64 201
rect 65 200 66 201
rect 60 201 66 205
rect 60 205 61 206
rect 62 205 63 206
rect 63 205 64 206
rect 65 205 66 206
rect 400 500 401 501
rect 402 500 403 501
rect 403 500 404 501
rect 405 500 406 501
rect 400 501 406 505
rect 400 505 401 506
rect 402 505 403 506
rect 403 505 404 506
rect 405 505 406 506
rect 160 0 161 1
rect 162 0 163 1
rect 163 0 164 1
rect 165 0 166 1
rect 160 1 166 5
rect 160 5 161 6
rect 162 5 163 6
rect 163 5 164 6
rect 165 5 166 6
rect 280 80 281 81
rect 282 80 283 81
rect 283 80 284 81
rect 285 80 286 81
rect 280 81 286 85
rect 280 85 281 86
rect 282 85 283 86
rect 283 85 284 86
rect 285 85 286 86
rect 40 180 41 181
rect 42 180 43 181
rect 43 180 44 181
rect 45 180 46 181
rect 40 181 46 185
rect 40 185 41 186
rect 42 185 43 186
rect 43 185 44 186
rect 45 185 46 186
rect 660 180 661 181
rect 662 180 663 181
rect 663 180 664 181
rect 665 180 666 181
rect 660 181 666 185
rect 660 185 661 186
rect 662 185 663 186
rect 663 185 664 186
rect 665 185 666 186
rect 340 260 341 261
rect 342 260 343 261
rect 343 260 344 261
rect 345 260 346 261
rect 340 261 346 265
rect 340 265 341 266
rect 342 265 343 266
rect 343 265 344 266
rect 345 265 346 266
rect 540 360 541 361
rect 542 360 543 361
rect 543 360 544 361
rect 545 360 546 361
rect 540 361 546 365
rect 540 365 541 366
rect 542 365 543 366
rect 543 365 544 366
rect 545 365 546 366
rect 80 80 81 81
rect 82 80 83 81
rect 83 80 84 81
rect 85 80 86 81
rect 80 81 86 85
rect 80 85 81 86
rect 82 85 83 86
rect 83 85 84 86
rect 85 85 86 86
rect 140 620 141 621
rect 142 620 143 621
rect 143 620 144 621
rect 145 620 146 621
rect 140 621 146 625
rect 140 625 141 626
rect 142 625 143 626
rect 143 625 144 626
rect 145 625 146 626
rect 480 80 481 81
rect 482 80 483 81
rect 483 80 484 81
rect 485 80 486 81
rect 480 81 486 85
rect 480 85 481 86
rect 482 85 483 86
rect 483 85 484 86
rect 485 85 486 86
rect 160 80 161 81
rect 162 80 163 81
rect 163 80 164 81
rect 165 80 166 81
rect 160 81 166 85
rect 160 85 161 86
rect 162 85 163 86
rect 163 85 164 86
rect 165 85 166 86
rect 260 660 261 661
rect 262 660 263 661
rect 263 660 264 661
rect 265 660 266 661
rect 260 661 266 665
rect 260 665 261 666
rect 262 665 263 666
rect 263 665 264 666
rect 265 665 266 666
rect 620 440 621 441
rect 622 440 623 441
rect 623 440 624 441
rect 625 440 626 441
rect 620 441 626 445
rect 620 445 621 446
rect 622 445 623 446
rect 623 445 624 446
rect 625 445 626 446
rect 100 280 101 281
rect 102 280 103 281
rect 103 280 104 281
rect 105 280 106 281
rect 100 281 106 285
rect 100 285 101 286
rect 102 285 103 286
rect 103 285 104 286
rect 105 285 106 286
rect 260 320 261 321
rect 262 320 263 321
rect 263 320 264 321
rect 265 320 266 321
rect 260 321 266 325
rect 260 325 261 326
rect 262 325 263 326
rect 263 325 264 326
rect 265 325 266 326
rect 500 400 501 401
rect 502 400 503 401
rect 503 400 504 401
rect 505 400 506 401
rect 500 401 506 405
rect 500 405 501 406
rect 502 405 503 406
rect 503 405 504 406
rect 505 405 506 406
rect 180 500 181 501
rect 182 500 183 501
rect 183 500 184 501
rect 185 500 186 501
rect 180 501 186 505
rect 180 505 181 506
rect 182 505 183 506
rect 183 505 184 506
rect 185 505 186 506
rect 260 520 261 521
rect 262 520 263 521
rect 263 520 264 521
rect 265 520 266 521
rect 260 521 266 525
rect 260 525 261 526
rect 262 525 263 526
rect 263 525 264 526
rect 265 525 266 526
rect 120 460 121 461
rect 122 460 123 461
rect 123 460 124 461
rect 125 460 126 461
rect 120 461 126 465
rect 120 465 121 466
rect 122 465 123 466
rect 123 465 124 466
rect 125 465 126 466
rect 620 360 621 361
rect 622 360 623 361
rect 623 360 624 361
rect 625 360 626 361
rect 620 361 626 365
rect 620 365 621 366
rect 622 365 623 366
rect 623 365 624 366
rect 625 365 626 366
rect 620 380 621 381
rect 622 380 623 381
rect 623 380 624 381
rect 625 380 626 381
rect 620 381 626 385
rect 620 385 621 386
rect 622 385 623 386
rect 623 385 624 386
rect 625 385 626 386
rect 540 180 541 181
rect 542 180 543 181
rect 543 180 544 181
rect 545 180 546 181
rect 540 181 546 185
rect 540 185 541 186
rect 542 185 543 186
rect 543 185 544 186
rect 545 185 546 186
rect 180 80 181 81
rect 182 80 183 81
rect 183 80 184 81
rect 185 80 186 81
rect 180 81 186 85
rect 180 85 181 86
rect 182 85 183 86
rect 183 85 184 86
rect 185 85 186 86
rect 200 500 201 501
rect 202 500 203 501
rect 203 500 204 501
rect 205 500 206 501
rect 200 501 206 505
rect 200 505 201 506
rect 202 505 203 506
rect 203 505 204 506
rect 205 505 206 506
rect 540 100 541 101
rect 542 100 543 101
rect 543 100 544 101
rect 545 100 546 101
rect 540 101 546 105
rect 540 105 541 106
rect 542 105 543 106
rect 543 105 544 106
rect 545 105 546 106
rect 260 200 261 201
rect 262 200 263 201
rect 263 200 264 201
rect 265 200 266 201
rect 260 201 266 205
rect 260 205 261 206
rect 262 205 263 206
rect 263 205 264 206
rect 265 205 266 206
rect 540 80 541 81
rect 542 80 543 81
rect 543 80 544 81
rect 545 80 546 81
rect 540 81 546 85
rect 540 85 541 86
rect 542 85 543 86
rect 543 85 544 86
rect 545 85 546 86
rect 220 340 221 341
rect 222 340 223 341
rect 223 340 224 341
rect 225 340 226 341
rect 220 341 226 345
rect 220 345 221 346
rect 222 345 223 346
rect 223 345 224 346
rect 225 345 226 346
rect 580 360 581 361
rect 582 360 583 361
rect 583 360 584 361
rect 585 360 586 361
rect 580 361 586 365
rect 580 365 581 366
rect 582 365 583 366
rect 583 365 584 366
rect 585 365 586 366
rect 600 200 601 201
rect 602 200 603 201
rect 603 200 604 201
rect 605 200 606 201
rect 600 201 606 205
rect 600 205 601 206
rect 602 205 603 206
rect 603 205 604 206
rect 605 205 606 206
rect 100 160 101 161
rect 102 160 103 161
rect 103 160 104 161
rect 105 160 106 161
rect 100 161 106 165
rect 100 165 101 166
rect 102 165 103 166
rect 103 165 104 166
rect 105 165 106 166
rect 40 540 41 541
rect 42 540 43 541
rect 43 540 44 541
rect 45 540 46 541
rect 40 541 46 545
rect 40 545 41 546
rect 42 545 43 546
rect 43 545 44 546
rect 45 545 46 546
rect 580 440 581 441
rect 582 440 583 441
rect 583 440 584 441
rect 585 440 586 441
rect 580 441 586 445
rect 580 445 581 446
rect 582 445 583 446
rect 583 445 584 446
rect 585 445 586 446
rect 80 520 81 521
rect 82 520 83 521
rect 83 520 84 521
rect 85 520 86 521
rect 80 521 86 525
rect 80 525 81 526
rect 82 525 83 526
rect 83 525 84 526
rect 85 525 86 526
rect 140 280 141 281
rect 142 280 143 281
rect 143 280 144 281
rect 145 280 146 281
rect 140 281 146 285
rect 140 285 141 286
rect 142 285 143 286
rect 143 285 144 286
rect 145 285 146 286
rect 240 600 241 601
rect 242 600 243 601
rect 243 600 244 601
rect 245 600 246 601
rect 240 601 246 605
rect 240 605 241 606
rect 242 605 243 606
rect 243 605 244 606
rect 245 605 246 606
rect 280 260 281 261
rect 282 260 283 261
rect 283 260 284 261
rect 285 260 286 261
rect 280 261 286 265
rect 280 265 281 266
rect 282 265 283 266
rect 283 265 284 266
rect 285 265 286 266
rect 160 540 161 541
rect 162 540 163 541
rect 163 540 164 541
rect 165 540 166 541
rect 160 541 166 545
rect 160 545 161 546
rect 162 545 163 546
rect 163 545 164 546
rect 165 545 166 546
rect 360 440 361 441
rect 362 440 363 441
rect 363 440 364 441
rect 365 440 366 441
rect 360 441 366 445
rect 360 445 361 446
rect 362 445 363 446
rect 363 445 364 446
rect 365 445 366 446
rect 220 80 221 81
rect 222 80 223 81
rect 223 80 224 81
rect 225 80 226 81
rect 220 81 226 85
rect 220 85 221 86
rect 222 85 223 86
rect 223 85 224 86
rect 225 85 226 86
rect 400 660 401 661
rect 402 660 403 661
rect 403 660 404 661
rect 405 660 406 661
rect 400 661 406 665
rect 400 665 401 666
rect 402 665 403 666
rect 403 665 404 666
rect 405 665 406 666
rect 0 440 1 441
rect 2 440 3 441
rect 3 440 4 441
rect 5 440 6 441
rect 0 441 6 445
rect 0 445 1 446
rect 2 445 3 446
rect 3 445 4 446
rect 5 445 6 446
rect 60 460 61 461
rect 62 460 63 461
rect 63 460 64 461
rect 65 460 66 461
rect 60 461 66 465
rect 60 465 61 466
rect 62 465 63 466
rect 63 465 64 466
rect 65 465 66 466
rect 540 480 541 481
rect 542 480 543 481
rect 543 480 544 481
rect 545 480 546 481
rect 540 481 546 485
rect 540 485 541 486
rect 542 485 543 486
rect 543 485 544 486
rect 545 485 546 486
rect 160 620 161 621
rect 162 620 163 621
rect 163 620 164 621
rect 165 620 166 621
rect 160 621 166 625
rect 160 625 161 626
rect 162 625 163 626
rect 163 625 164 626
rect 165 625 166 626
rect 180 580 181 581
rect 182 580 183 581
rect 183 580 184 581
rect 185 580 186 581
rect 180 581 186 585
rect 180 585 181 586
rect 182 585 183 586
rect 183 585 184 586
rect 185 585 186 586
rect 0 400 1 401
rect 2 400 3 401
rect 3 400 4 401
rect 5 400 6 401
rect 0 401 6 405
rect 0 405 1 406
rect 2 405 3 406
rect 3 405 4 406
rect 5 405 6 406
rect 280 140 281 141
rect 282 140 283 141
rect 283 140 284 141
rect 285 140 286 141
rect 280 141 286 145
rect 280 145 281 146
rect 282 145 283 146
rect 283 145 284 146
rect 285 145 286 146
rect 460 280 461 281
rect 462 280 463 281
rect 463 280 464 281
rect 465 280 466 281
rect 460 281 466 285
rect 460 285 461 286
rect 462 285 463 286
rect 463 285 464 286
rect 465 285 466 286
rect 420 60 421 61
rect 422 60 423 61
rect 423 60 424 61
rect 425 60 426 61
rect 420 61 426 65
rect 420 65 421 66
rect 422 65 423 66
rect 423 65 424 66
rect 425 65 426 66
rect 100 300 101 301
rect 102 300 103 301
rect 103 300 104 301
rect 105 300 106 301
rect 100 301 106 305
rect 100 305 101 306
rect 102 305 103 306
rect 103 305 104 306
rect 105 305 106 306
rect 360 120 361 121
rect 362 120 363 121
rect 363 120 364 121
rect 365 120 366 121
rect 360 121 366 125
rect 360 125 361 126
rect 362 125 363 126
rect 363 125 364 126
rect 365 125 366 126
rect 0 140 1 141
rect 2 140 3 141
rect 3 140 4 141
rect 5 140 6 141
rect 0 141 6 145
rect 0 145 1 146
rect 2 145 3 146
rect 3 145 4 146
rect 5 145 6 146
rect 500 200 501 201
rect 502 200 503 201
rect 503 200 504 201
rect 505 200 506 201
rect 500 201 506 205
rect 500 205 501 206
rect 502 205 503 206
rect 503 205 504 206
rect 505 205 506 206
rect 60 260 61 261
rect 62 260 63 261
rect 63 260 64 261
rect 65 260 66 261
rect 60 261 66 265
rect 60 265 61 266
rect 62 265 63 266
rect 63 265 64 266
rect 65 265 66 266
rect 400 260 401 261
rect 402 260 403 261
rect 403 260 404 261
rect 405 260 406 261
rect 400 261 406 265
rect 400 265 401 266
rect 402 265 403 266
rect 403 265 404 266
rect 405 265 406 266
rect 580 380 581 381
rect 582 380 583 381
rect 583 380 584 381
rect 585 380 586 381
rect 580 381 586 385
rect 580 385 581 386
rect 582 385 583 386
rect 583 385 584 386
rect 585 385 586 386
rect 100 600 101 601
rect 102 600 103 601
rect 103 600 104 601
rect 105 600 106 601
rect 100 601 106 605
rect 100 605 101 606
rect 102 605 103 606
rect 103 605 104 606
rect 105 605 106 606
rect 600 320 601 321
rect 602 320 603 321
rect 603 320 604 321
rect 605 320 606 321
rect 600 321 606 325
rect 600 325 601 326
rect 602 325 603 326
rect 603 325 604 326
rect 605 325 606 326
rect 160 480 161 481
rect 162 480 163 481
rect 163 480 164 481
rect 165 480 166 481
rect 160 481 166 485
rect 160 485 161 486
rect 162 485 163 486
rect 163 485 164 486
rect 165 485 166 486
rect 140 420 141 421
rect 142 420 143 421
rect 143 420 144 421
rect 145 420 146 421
rect 140 421 146 425
rect 140 425 141 426
rect 142 425 143 426
rect 143 425 144 426
rect 145 425 146 426
rect 260 360 261 361
rect 262 360 263 361
rect 263 360 264 361
rect 265 360 266 361
rect 260 361 266 365
rect 260 365 261 366
rect 262 365 263 366
rect 263 365 264 366
rect 265 365 266 366
rect 120 360 121 361
rect 122 360 123 361
rect 123 360 124 361
rect 125 360 126 361
rect 120 361 126 365
rect 120 365 121 366
rect 122 365 123 366
rect 123 365 124 366
rect 125 365 126 366
rect 340 280 341 281
rect 342 280 343 281
rect 343 280 344 281
rect 345 280 346 281
rect 340 281 346 285
rect 340 285 341 286
rect 342 285 343 286
rect 343 285 344 286
rect 345 285 346 286
rect 100 580 101 581
rect 102 580 103 581
rect 103 580 104 581
rect 105 580 106 581
rect 100 581 106 585
rect 100 585 101 586
rect 102 585 103 586
rect 103 585 104 586
rect 105 585 106 586
rect 100 340 101 341
rect 102 340 103 341
rect 103 340 104 341
rect 105 340 106 341
rect 100 341 106 345
rect 100 345 101 346
rect 102 345 103 346
rect 103 345 104 346
rect 105 345 106 346
rect 520 460 521 461
rect 522 460 523 461
rect 523 460 524 461
rect 525 460 526 461
rect 520 461 526 465
rect 520 465 521 466
rect 522 465 523 466
rect 523 465 524 466
rect 525 465 526 466
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect 620 240 621 241
rect 622 240 623 241
rect 623 240 624 241
rect 625 240 626 241
rect 620 241 626 245
rect 620 245 621 246
rect 622 245 623 246
rect 623 245 624 246
rect 625 245 626 246
rect 120 220 121 221
rect 122 220 123 221
rect 123 220 124 221
rect 125 220 126 221
rect 120 221 126 225
rect 120 225 121 226
rect 122 225 123 226
rect 123 225 124 226
rect 125 225 126 226
rect 360 20 361 21
rect 362 20 363 21
rect 363 20 364 21
rect 365 20 366 21
rect 360 21 366 25
rect 360 25 361 26
rect 362 25 363 26
rect 363 25 364 26
rect 365 25 366 26
rect 380 220 381 221
rect 382 220 383 221
rect 383 220 384 221
rect 385 220 386 221
rect 380 221 386 225
rect 380 225 381 226
rect 382 225 383 226
rect 383 225 384 226
rect 385 225 386 226
rect 100 60 101 61
rect 102 60 103 61
rect 103 60 104 61
rect 105 60 106 61
rect 100 61 106 65
rect 100 65 101 66
rect 102 65 103 66
rect 103 65 104 66
rect 105 65 106 66
rect 640 400 641 401
rect 642 400 643 401
rect 643 400 644 401
rect 645 400 646 401
rect 640 401 646 405
rect 640 405 641 406
rect 642 405 643 406
rect 643 405 644 406
rect 645 405 646 406
rect 40 360 41 361
rect 42 360 43 361
rect 43 360 44 361
rect 45 360 46 361
rect 40 361 46 365
rect 40 365 41 366
rect 42 365 43 366
rect 43 365 44 366
rect 45 365 46 366
rect 500 520 501 521
rect 502 520 503 521
rect 503 520 504 521
rect 505 520 506 521
rect 500 521 506 525
rect 500 525 501 526
rect 502 525 503 526
rect 503 525 504 526
rect 505 525 506 526
rect 240 160 241 161
rect 242 160 243 161
rect 243 160 244 161
rect 245 160 246 161
rect 240 161 246 165
rect 240 165 241 166
rect 242 165 243 166
rect 243 165 244 166
rect 245 165 246 166
rect 620 220 621 221
rect 622 220 623 221
rect 623 220 624 221
rect 625 220 626 221
rect 620 221 626 225
rect 620 225 621 226
rect 622 225 623 226
rect 623 225 624 226
rect 625 225 626 226
rect 400 320 401 321
rect 402 320 403 321
rect 403 320 404 321
rect 405 320 406 321
rect 400 321 406 325
rect 400 325 401 326
rect 402 325 403 326
rect 403 325 404 326
rect 405 325 406 326
rect 360 60 361 61
rect 362 60 363 61
rect 363 60 364 61
rect 365 60 366 61
rect 360 61 366 65
rect 360 65 361 66
rect 362 65 363 66
rect 363 65 364 66
rect 365 65 366 66
rect 600 460 601 461
rect 602 460 603 461
rect 603 460 604 461
rect 605 460 606 461
rect 600 461 606 465
rect 600 465 601 466
rect 602 465 603 466
rect 603 465 604 466
rect 605 465 606 466
rect 400 20 401 21
rect 402 20 403 21
rect 403 20 404 21
rect 405 20 406 21
rect 400 21 406 25
rect 400 25 401 26
rect 402 25 403 26
rect 403 25 404 26
rect 405 25 406 26
rect 580 220 581 221
rect 582 220 583 221
rect 583 220 584 221
rect 585 220 586 221
rect 580 221 586 225
rect 580 225 581 226
rect 582 225 583 226
rect 583 225 584 226
rect 585 225 586 226
rect 480 0 481 1
rect 482 0 483 1
rect 483 0 484 1
rect 485 0 486 1
rect 480 1 486 5
rect 480 5 481 6
rect 482 5 483 6
rect 483 5 484 6
rect 485 5 486 6
rect 520 120 521 121
rect 522 120 523 121
rect 523 120 524 121
rect 525 120 526 121
rect 520 121 526 125
rect 520 125 521 126
rect 522 125 523 126
rect 523 125 524 126
rect 525 125 526 126
rect 600 420 601 421
rect 602 420 603 421
rect 603 420 604 421
rect 605 420 606 421
rect 600 421 606 425
rect 600 425 601 426
rect 602 425 603 426
rect 603 425 604 426
rect 605 425 606 426
rect 400 400 401 401
rect 402 400 403 401
rect 403 400 404 401
rect 405 400 406 401
rect 400 401 406 405
rect 400 405 401 406
rect 402 405 403 406
rect 403 405 404 406
rect 405 405 406 406
rect 340 40 341 41
rect 342 40 343 41
rect 343 40 344 41
rect 345 40 346 41
rect 340 41 346 45
rect 340 45 341 46
rect 342 45 343 46
rect 343 45 344 46
rect 345 45 346 46
rect 320 360 321 361
rect 322 360 323 361
rect 323 360 324 361
rect 325 360 326 361
rect 320 361 326 365
rect 320 365 321 366
rect 322 365 323 366
rect 323 365 324 366
rect 325 365 326 366
rect 160 40 161 41
rect 162 40 163 41
rect 163 40 164 41
rect 165 40 166 41
rect 160 41 166 45
rect 160 45 161 46
rect 162 45 163 46
rect 163 45 164 46
rect 165 45 166 46
rect 40 160 41 161
rect 42 160 43 161
rect 43 160 44 161
rect 45 160 46 161
rect 40 161 46 165
rect 40 165 41 166
rect 42 165 43 166
rect 43 165 44 166
rect 45 165 46 166
rect 120 180 121 181
rect 122 180 123 181
rect 123 180 124 181
rect 125 180 126 181
rect 120 181 126 185
rect 120 185 121 186
rect 122 185 123 186
rect 123 185 124 186
rect 125 185 126 186
rect 280 620 281 621
rect 282 620 283 621
rect 283 620 284 621
rect 285 620 286 621
rect 280 621 286 625
rect 280 625 281 626
rect 282 625 283 626
rect 283 625 284 626
rect 285 625 286 626
rect 180 600 181 601
rect 182 600 183 601
rect 183 600 184 601
rect 185 600 186 601
rect 180 601 186 605
rect 180 605 181 606
rect 182 605 183 606
rect 183 605 184 606
rect 185 605 186 606
rect 580 120 581 121
rect 582 120 583 121
rect 583 120 584 121
rect 585 120 586 121
rect 580 121 586 125
rect 580 125 581 126
rect 582 125 583 126
rect 583 125 584 126
rect 585 125 586 126
rect 300 620 301 621
rect 302 620 303 621
rect 303 620 304 621
rect 305 620 306 621
rect 300 621 306 625
rect 300 625 301 626
rect 302 625 303 626
rect 303 625 304 626
rect 305 625 306 626
rect 80 380 81 381
rect 82 380 83 381
rect 83 380 84 381
rect 85 380 86 381
rect 80 381 86 385
rect 80 385 81 386
rect 82 385 83 386
rect 83 385 84 386
rect 85 385 86 386
rect 640 420 641 421
rect 642 420 643 421
rect 643 420 644 421
rect 645 420 646 421
rect 640 421 646 425
rect 640 425 641 426
rect 642 425 643 426
rect 643 425 644 426
rect 645 425 646 426
rect 320 560 321 561
rect 322 560 323 561
rect 323 560 324 561
rect 325 560 326 561
rect 320 561 326 565
rect 320 565 321 566
rect 322 565 323 566
rect 323 565 324 566
rect 325 565 326 566
rect 420 340 421 341
rect 422 340 423 341
rect 423 340 424 341
rect 425 340 426 341
rect 420 341 426 345
rect 420 345 421 346
rect 422 345 423 346
rect 423 345 424 346
rect 425 345 426 346
rect 60 480 61 481
rect 62 480 63 481
rect 63 480 64 481
rect 65 480 66 481
rect 60 481 66 485
rect 60 485 61 486
rect 62 485 63 486
rect 63 485 64 486
rect 65 485 66 486
rect 660 400 661 401
rect 662 400 663 401
rect 663 400 664 401
rect 665 400 666 401
rect 660 401 666 405
rect 660 405 661 406
rect 662 405 663 406
rect 663 405 664 406
rect 665 405 666 406
rect 220 20 221 21
rect 222 20 223 21
rect 223 20 224 21
rect 225 20 226 21
rect 220 21 226 25
rect 220 25 221 26
rect 222 25 223 26
rect 223 25 224 26
rect 225 25 226 26
rect 0 120 1 121
rect 2 120 3 121
rect 3 120 4 121
rect 5 120 6 121
rect 0 121 6 125
rect 0 125 1 126
rect 2 125 3 126
rect 3 125 4 126
rect 5 125 6 126
rect 520 400 521 401
rect 522 400 523 401
rect 523 400 524 401
rect 525 400 526 401
rect 520 401 526 405
rect 520 405 521 406
rect 522 405 523 406
rect 523 405 524 406
rect 525 405 526 406
rect 20 480 21 481
rect 22 480 23 481
rect 23 480 24 481
rect 25 480 26 481
rect 20 481 26 485
rect 20 485 21 486
rect 22 485 23 486
rect 23 485 24 486
rect 25 485 26 486
rect 180 340 181 341
rect 182 340 183 341
rect 183 340 184 341
rect 185 340 186 341
rect 180 341 186 345
rect 180 345 181 346
rect 182 345 183 346
rect 183 345 184 346
rect 185 345 186 346
rect 560 480 561 481
rect 562 480 563 481
rect 563 480 564 481
rect 565 480 566 481
rect 560 481 566 485
rect 560 485 561 486
rect 562 485 563 486
rect 563 485 564 486
rect 565 485 566 486
rect 420 180 421 181
rect 422 180 423 181
rect 423 180 424 181
rect 425 180 426 181
rect 420 181 426 185
rect 420 185 421 186
rect 422 185 423 186
rect 423 185 424 186
rect 425 185 426 186
rect 280 200 281 201
rect 282 200 283 201
rect 283 200 284 201
rect 285 200 286 201
rect 280 201 286 205
rect 280 205 281 206
rect 282 205 283 206
rect 283 205 284 206
rect 285 205 286 206
rect 480 40 481 41
rect 482 40 483 41
rect 483 40 484 41
rect 485 40 486 41
rect 480 41 486 45
rect 480 45 481 46
rect 482 45 483 46
rect 483 45 484 46
rect 485 45 486 46
rect 60 220 61 221
rect 62 220 63 221
rect 63 220 64 221
rect 65 220 66 221
rect 60 221 66 225
rect 60 225 61 226
rect 62 225 63 226
rect 63 225 64 226
rect 65 225 66 226
rect 140 600 141 601
rect 142 600 143 601
rect 143 600 144 601
rect 145 600 146 601
rect 140 601 146 605
rect 140 605 141 606
rect 142 605 143 606
rect 143 605 144 606
rect 145 605 146 606
rect 140 560 141 561
rect 142 560 143 561
rect 143 560 144 561
rect 145 560 146 561
rect 140 561 146 565
rect 140 565 141 566
rect 142 565 143 566
rect 143 565 144 566
rect 145 565 146 566
rect 100 120 101 121
rect 102 120 103 121
rect 103 120 104 121
rect 105 120 106 121
rect 100 121 106 125
rect 100 125 101 126
rect 102 125 103 126
rect 103 125 104 126
rect 105 125 106 126
rect 480 380 481 381
rect 482 380 483 381
rect 483 380 484 381
rect 485 380 486 381
rect 480 381 486 385
rect 480 385 481 386
rect 482 385 483 386
rect 483 385 484 386
rect 485 385 486 386
rect 660 420 661 421
rect 662 420 663 421
rect 663 420 664 421
rect 665 420 666 421
rect 660 421 666 425
rect 660 425 661 426
rect 662 425 663 426
rect 663 425 664 426
rect 665 425 666 426
rect 160 60 161 61
rect 162 60 163 61
rect 163 60 164 61
rect 165 60 166 61
rect 160 61 166 65
rect 160 65 161 66
rect 162 65 163 66
rect 163 65 164 66
rect 165 65 166 66
rect 0 520 1 521
rect 2 520 3 521
rect 3 520 4 521
rect 5 520 6 521
rect 0 521 6 525
rect 0 525 1 526
rect 2 525 3 526
rect 3 525 4 526
rect 5 525 6 526
rect 560 360 561 361
rect 562 360 563 361
rect 563 360 564 361
rect 565 360 566 361
rect 560 361 566 365
rect 560 365 561 366
rect 562 365 563 366
rect 563 365 564 366
rect 565 365 566 366
rect 40 120 41 121
rect 42 120 43 121
rect 43 120 44 121
rect 45 120 46 121
rect 40 121 46 125
rect 40 125 41 126
rect 42 125 43 126
rect 43 125 44 126
rect 45 125 46 126
rect 140 300 141 301
rect 142 300 143 301
rect 143 300 144 301
rect 145 300 146 301
rect 140 301 146 305
rect 140 305 141 306
rect 142 305 143 306
rect 143 305 144 306
rect 145 305 146 306
rect 0 420 1 421
rect 2 420 3 421
rect 3 420 4 421
rect 5 420 6 421
rect 0 421 6 425
rect 0 425 1 426
rect 2 425 3 426
rect 3 425 4 426
rect 5 425 6 426
rect 80 220 81 221
rect 82 220 83 221
rect 83 220 84 221
rect 85 220 86 221
rect 80 221 86 225
rect 80 225 81 226
rect 82 225 83 226
rect 83 225 84 226
rect 85 225 86 226
rect 20 120 21 121
rect 22 120 23 121
rect 23 120 24 121
rect 25 120 26 121
rect 20 121 26 125
rect 20 125 21 126
rect 22 125 23 126
rect 23 125 24 126
rect 25 125 26 126
rect 260 640 261 641
rect 262 640 263 641
rect 263 640 264 641
rect 265 640 266 641
rect 260 641 266 645
rect 260 645 261 646
rect 262 645 263 646
rect 263 645 264 646
rect 265 645 266 646
rect 420 480 421 481
rect 422 480 423 481
rect 423 480 424 481
rect 425 480 426 481
rect 420 481 426 485
rect 420 485 421 486
rect 422 485 423 486
rect 423 485 424 486
rect 425 485 426 486
rect 380 40 381 41
rect 382 40 383 41
rect 383 40 384 41
rect 385 40 386 41
rect 380 41 386 45
rect 380 45 381 46
rect 382 45 383 46
rect 383 45 384 46
rect 385 45 386 46
rect 200 660 201 661
rect 202 660 203 661
rect 203 660 204 661
rect 205 660 206 661
rect 200 661 206 665
rect 200 665 201 666
rect 202 665 203 666
rect 203 665 204 666
rect 205 665 206 666
rect 440 500 441 501
rect 442 500 443 501
rect 443 500 444 501
rect 445 500 446 501
rect 440 501 446 505
rect 440 505 441 506
rect 442 505 443 506
rect 443 505 444 506
rect 445 505 446 506
rect 460 120 461 121
rect 462 120 463 121
rect 463 120 464 121
rect 465 120 466 121
rect 460 121 466 125
rect 460 125 461 126
rect 462 125 463 126
rect 463 125 464 126
rect 465 125 466 126
rect 160 200 161 201
rect 162 200 163 201
rect 163 200 164 201
rect 165 200 166 201
rect 160 201 166 205
rect 160 205 161 206
rect 162 205 163 206
rect 163 205 164 206
rect 165 205 166 206
rect 240 40 241 41
rect 242 40 243 41
rect 243 40 244 41
rect 245 40 246 41
rect 240 41 246 45
rect 240 45 241 46
rect 242 45 243 46
rect 243 45 244 46
rect 245 45 246 46
rect 300 520 301 521
rect 302 520 303 521
rect 303 520 304 521
rect 305 520 306 521
rect 300 521 306 525
rect 300 525 301 526
rect 302 525 303 526
rect 303 525 304 526
rect 305 525 306 526
rect 500 600 501 601
rect 502 600 503 601
rect 503 600 504 601
rect 505 600 506 601
rect 500 601 506 605
rect 500 605 501 606
rect 502 605 503 606
rect 503 605 504 606
rect 505 605 506 606
rect 320 260 321 261
rect 322 260 323 261
rect 323 260 324 261
rect 325 260 326 261
rect 320 261 326 265
rect 320 265 321 266
rect 322 265 323 266
rect 323 265 324 266
rect 325 265 326 266
rect 600 360 601 361
rect 602 360 603 361
rect 603 360 604 361
rect 605 360 606 361
rect 600 361 606 365
rect 600 365 601 366
rect 602 365 603 366
rect 603 365 604 366
rect 605 365 606 366
rect 580 260 581 261
rect 582 260 583 261
rect 583 260 584 261
rect 585 260 586 261
rect 580 261 586 265
rect 580 265 581 266
rect 582 265 583 266
rect 583 265 584 266
rect 585 265 586 266
rect 320 660 321 661
rect 322 660 323 661
rect 323 660 324 661
rect 325 660 326 661
rect 320 661 326 665
rect 320 665 321 666
rect 322 665 323 666
rect 323 665 324 666
rect 325 665 326 666
rect 560 160 561 161
rect 562 160 563 161
rect 563 160 564 161
rect 565 160 566 161
rect 560 161 566 165
rect 560 165 561 166
rect 562 165 563 166
rect 563 165 564 166
rect 565 165 566 166
rect 480 280 481 281
rect 482 280 483 281
rect 483 280 484 281
rect 485 280 486 281
rect 480 281 486 285
rect 480 285 481 286
rect 482 285 483 286
rect 483 285 484 286
rect 485 285 486 286
rect 460 540 461 541
rect 462 540 463 541
rect 463 540 464 541
rect 465 540 466 541
rect 460 541 466 545
rect 460 545 461 546
rect 462 545 463 546
rect 463 545 464 546
rect 465 545 466 546
rect 0 300 1 301
rect 2 300 3 301
rect 3 300 4 301
rect 5 300 6 301
rect 0 301 6 305
rect 0 305 1 306
rect 2 305 3 306
rect 3 305 4 306
rect 5 305 6 306
rect 60 280 61 281
rect 62 280 63 281
rect 63 280 64 281
rect 65 280 66 281
rect 60 281 66 285
rect 60 285 61 286
rect 62 285 63 286
rect 63 285 64 286
rect 65 285 66 286
rect 380 320 381 321
rect 382 320 383 321
rect 383 320 384 321
rect 385 320 386 321
rect 380 321 386 325
rect 380 325 381 326
rect 382 325 383 326
rect 383 325 384 326
rect 385 325 386 326
rect 120 560 121 561
rect 122 560 123 561
rect 123 560 124 561
rect 125 560 126 561
rect 120 561 126 565
rect 120 565 121 566
rect 122 565 123 566
rect 123 565 124 566
rect 125 565 126 566
rect 640 200 641 201
rect 642 200 643 201
rect 643 200 644 201
rect 645 200 646 201
rect 640 201 646 205
rect 640 205 641 206
rect 642 205 643 206
rect 643 205 644 206
rect 645 205 646 206
rect 180 420 181 421
rect 182 420 183 421
rect 183 420 184 421
rect 185 420 186 421
rect 180 421 186 425
rect 180 425 181 426
rect 182 425 183 426
rect 183 425 184 426
rect 185 425 186 426
rect 380 640 381 641
rect 382 640 383 641
rect 383 640 384 641
rect 385 640 386 641
rect 380 641 386 645
rect 380 645 381 646
rect 382 645 383 646
rect 383 645 384 646
rect 385 645 386 646
rect 240 400 241 401
rect 242 400 243 401
rect 243 400 244 401
rect 245 400 246 401
rect 240 401 246 405
rect 240 405 241 406
rect 242 405 243 406
rect 243 405 244 406
rect 245 405 246 406
rect 220 400 221 401
rect 222 400 223 401
rect 223 400 224 401
rect 225 400 226 401
rect 220 401 226 405
rect 220 405 221 406
rect 222 405 223 406
rect 223 405 224 406
rect 225 405 226 406
rect 200 280 201 281
rect 202 280 203 281
rect 203 280 204 281
rect 205 280 206 281
rect 200 281 206 285
rect 200 285 201 286
rect 202 285 203 286
rect 203 285 204 286
rect 205 285 206 286
rect 560 500 561 501
rect 562 500 563 501
rect 563 500 564 501
rect 565 500 566 501
rect 560 501 566 505
rect 560 505 561 506
rect 562 505 563 506
rect 563 505 564 506
rect 565 505 566 506
rect 20 420 21 421
rect 22 420 23 421
rect 23 420 24 421
rect 25 420 26 421
rect 20 421 26 425
rect 20 425 21 426
rect 22 425 23 426
rect 23 425 24 426
rect 25 425 26 426
rect 460 440 461 441
rect 462 440 463 441
rect 463 440 464 441
rect 465 440 466 441
rect 460 441 466 445
rect 460 445 461 446
rect 462 445 463 446
rect 463 445 464 446
rect 465 445 466 446
rect 520 320 521 321
rect 522 320 523 321
rect 523 320 524 321
rect 525 320 526 321
rect 520 321 526 325
rect 520 325 521 326
rect 522 325 523 326
rect 523 325 524 326
rect 525 325 526 326
rect 460 300 461 301
rect 462 300 463 301
rect 463 300 464 301
rect 465 300 466 301
rect 460 301 466 305
rect 460 305 461 306
rect 462 305 463 306
rect 463 305 464 306
rect 465 305 466 306
rect 280 360 281 361
rect 282 360 283 361
rect 283 360 284 361
rect 285 360 286 361
rect 280 361 286 365
rect 280 365 281 366
rect 282 365 283 366
rect 283 365 284 366
rect 285 365 286 366
rect 240 20 241 21
rect 242 20 243 21
rect 243 20 244 21
rect 245 20 246 21
rect 240 21 246 25
rect 240 25 241 26
rect 242 25 243 26
rect 243 25 244 26
rect 245 25 246 26
rect 260 280 261 281
rect 262 280 263 281
rect 263 280 264 281
rect 265 280 266 281
rect 260 281 266 285
rect 260 285 261 286
rect 262 285 263 286
rect 263 285 264 286
rect 265 285 266 286
rect 240 100 241 101
rect 242 100 243 101
rect 243 100 244 101
rect 245 100 246 101
rect 240 101 246 105
rect 240 105 241 106
rect 242 105 243 106
rect 243 105 244 106
rect 245 105 246 106
rect 220 380 221 381
rect 222 380 223 381
rect 223 380 224 381
rect 225 380 226 381
rect 220 381 226 385
rect 220 385 221 386
rect 222 385 223 386
rect 223 385 224 386
rect 225 385 226 386
rect 560 240 561 241
rect 562 240 563 241
rect 563 240 564 241
rect 565 240 566 241
rect 560 241 566 245
rect 560 245 561 246
rect 562 245 563 246
rect 563 245 564 246
rect 565 245 566 246
rect 520 420 521 421
rect 522 420 523 421
rect 523 420 524 421
rect 525 420 526 421
rect 520 421 526 425
rect 520 425 521 426
rect 522 425 523 426
rect 523 425 524 426
rect 525 425 526 426
rect 440 620 441 621
rect 442 620 443 621
rect 443 620 444 621
rect 445 620 446 621
rect 440 621 446 625
rect 440 625 441 626
rect 442 625 443 626
rect 443 625 444 626
rect 445 625 446 626
rect 560 340 561 341
rect 562 340 563 341
rect 563 340 564 341
rect 565 340 566 341
rect 560 341 566 345
rect 560 345 561 346
rect 562 345 563 346
rect 563 345 564 346
rect 565 345 566 346
rect 180 640 181 641
rect 182 640 183 641
rect 183 640 184 641
rect 185 640 186 641
rect 180 641 186 645
rect 180 645 181 646
rect 182 645 183 646
rect 183 645 184 646
rect 185 645 186 646
rect 320 100 321 101
rect 322 100 323 101
rect 323 100 324 101
rect 325 100 326 101
rect 320 101 326 105
rect 320 105 321 106
rect 322 105 323 106
rect 323 105 324 106
rect 325 105 326 106
rect 440 280 441 281
rect 442 280 443 281
rect 443 280 444 281
rect 445 280 446 281
rect 440 281 446 285
rect 440 285 441 286
rect 442 285 443 286
rect 443 285 444 286
rect 445 285 446 286
rect 620 520 621 521
rect 622 520 623 521
rect 623 520 624 521
rect 625 520 626 521
rect 620 521 626 525
rect 620 525 621 526
rect 622 525 623 526
rect 623 525 624 526
rect 625 525 626 526
rect 180 400 181 401
rect 182 400 183 401
rect 183 400 184 401
rect 185 400 186 401
rect 180 401 186 405
rect 180 405 181 406
rect 182 405 183 406
rect 183 405 184 406
rect 185 405 186 406
rect 340 560 341 561
rect 342 560 343 561
rect 343 560 344 561
rect 345 560 346 561
rect 340 561 346 565
rect 340 565 341 566
rect 342 565 343 566
rect 343 565 344 566
rect 345 565 346 566
rect 300 420 301 421
rect 302 420 303 421
rect 303 420 304 421
rect 305 420 306 421
rect 300 421 306 425
rect 300 425 301 426
rect 302 425 303 426
rect 303 425 304 426
rect 305 425 306 426
rect 520 80 521 81
rect 522 80 523 81
rect 523 80 524 81
rect 525 80 526 81
rect 520 81 526 85
rect 520 85 521 86
rect 522 85 523 86
rect 523 85 524 86
rect 525 85 526 86
rect 520 500 521 501
rect 522 500 523 501
rect 523 500 524 501
rect 525 500 526 501
rect 520 501 526 505
rect 520 505 521 506
rect 522 505 523 506
rect 523 505 524 506
rect 525 505 526 506
rect 100 260 101 261
rect 102 260 103 261
rect 103 260 104 261
rect 105 260 106 261
rect 100 261 106 265
rect 100 265 101 266
rect 102 265 103 266
rect 103 265 104 266
rect 105 265 106 266
rect 120 260 121 261
rect 122 260 123 261
rect 123 260 124 261
rect 125 260 126 261
rect 120 261 126 265
rect 120 265 121 266
rect 122 265 123 266
rect 123 265 124 266
rect 125 265 126 266
rect 420 200 421 201
rect 422 200 423 201
rect 423 200 424 201
rect 425 200 426 201
rect 420 201 426 205
rect 420 205 421 206
rect 422 205 423 206
rect 423 205 424 206
rect 425 205 426 206
rect 140 320 141 321
rect 142 320 143 321
rect 143 320 144 321
rect 145 320 146 321
rect 140 321 146 325
rect 140 325 141 326
rect 142 325 143 326
rect 143 325 144 326
rect 145 325 146 326
rect 620 500 621 501
rect 622 500 623 501
rect 623 500 624 501
rect 625 500 626 501
rect 620 501 626 505
rect 620 505 621 506
rect 622 505 623 506
rect 623 505 624 506
rect 625 505 626 506
rect 160 340 161 341
rect 162 340 163 341
rect 163 340 164 341
rect 165 340 166 341
rect 160 341 166 345
rect 160 345 161 346
rect 162 345 163 346
rect 163 345 164 346
rect 165 345 166 346
rect 200 560 201 561
rect 202 560 203 561
rect 203 560 204 561
rect 205 560 206 561
rect 200 561 206 565
rect 200 565 201 566
rect 202 565 203 566
rect 203 565 204 566
rect 205 565 206 566
rect 200 220 201 221
rect 202 220 203 221
rect 203 220 204 221
rect 205 220 206 221
rect 200 221 206 225
rect 200 225 201 226
rect 202 225 203 226
rect 203 225 204 226
rect 205 225 206 226
rect 380 500 381 501
rect 382 500 383 501
rect 383 500 384 501
rect 385 500 386 501
rect 380 501 386 505
rect 380 505 381 506
rect 382 505 383 506
rect 383 505 384 506
rect 385 505 386 506
rect 520 60 521 61
rect 522 60 523 61
rect 523 60 524 61
rect 525 60 526 61
rect 520 61 526 65
rect 520 65 521 66
rect 522 65 523 66
rect 523 65 524 66
rect 525 65 526 66
rect 340 600 341 601
rect 342 600 343 601
rect 343 600 344 601
rect 345 600 346 601
rect 340 601 346 605
rect 340 605 341 606
rect 342 605 343 606
rect 343 605 344 606
rect 345 605 346 606
rect 380 160 381 161
rect 382 160 383 161
rect 383 160 384 161
rect 385 160 386 161
rect 380 161 386 165
rect 380 165 381 166
rect 382 165 383 166
rect 383 165 384 166
rect 385 165 386 166
rect 160 640 161 641
rect 162 640 163 641
rect 163 640 164 641
rect 165 640 166 641
rect 160 641 166 645
rect 160 645 161 646
rect 162 645 163 646
rect 163 645 164 646
rect 165 645 166 646
rect 220 520 221 521
rect 222 520 223 521
rect 223 520 224 521
rect 225 520 226 521
rect 220 521 226 525
rect 220 525 221 526
rect 222 525 223 526
rect 223 525 224 526
rect 225 525 226 526
rect 380 420 381 421
rect 382 420 383 421
rect 383 420 384 421
rect 385 420 386 421
rect 380 421 386 425
rect 380 425 381 426
rect 382 425 383 426
rect 383 425 384 426
rect 385 425 386 426
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect 500 440 501 441
rect 502 440 503 441
rect 503 440 504 441
rect 505 440 506 441
rect 500 441 506 445
rect 500 445 501 446
rect 502 445 503 446
rect 503 445 504 446
rect 505 445 506 446
rect 500 280 501 281
rect 502 280 503 281
rect 503 280 504 281
rect 505 280 506 281
rect 500 281 506 285
rect 500 285 501 286
rect 502 285 503 286
rect 503 285 504 286
rect 505 285 506 286
rect 640 340 641 341
rect 642 340 643 341
rect 643 340 644 341
rect 645 340 646 341
rect 640 341 646 345
rect 640 345 641 346
rect 642 345 643 346
rect 643 345 644 346
rect 645 345 646 346
rect 140 140 141 141
rect 142 140 143 141
rect 143 140 144 141
rect 145 140 146 141
rect 140 141 146 145
rect 140 145 141 146
rect 142 145 143 146
rect 143 145 144 146
rect 145 145 146 146
rect 360 640 361 641
rect 362 640 363 641
rect 363 640 364 641
rect 365 640 366 641
rect 360 641 366 645
rect 360 645 361 646
rect 362 645 363 646
rect 363 645 364 646
rect 365 645 366 646
rect 500 480 501 481
rect 502 480 503 481
rect 503 480 504 481
rect 505 480 506 481
rect 500 481 506 485
rect 500 485 501 486
rect 502 485 503 486
rect 503 485 504 486
rect 505 485 506 486
rect 380 280 381 281
rect 382 280 383 281
rect 383 280 384 281
rect 385 280 386 281
rect 380 281 386 285
rect 380 285 381 286
rect 382 285 383 286
rect 383 285 384 286
rect 385 285 386 286
rect 240 620 241 621
rect 242 620 243 621
rect 243 620 244 621
rect 245 620 246 621
rect 240 621 246 625
rect 240 625 241 626
rect 242 625 243 626
rect 243 625 244 626
rect 245 625 246 626
rect 260 560 261 561
rect 262 560 263 561
rect 263 560 264 561
rect 265 560 266 561
rect 260 561 266 565
rect 260 565 261 566
rect 262 565 263 566
rect 263 565 264 566
rect 265 565 266 566
rect 100 440 101 441
rect 102 440 103 441
rect 103 440 104 441
rect 105 440 106 441
rect 100 441 106 445
rect 100 445 101 446
rect 102 445 103 446
rect 103 445 104 446
rect 105 445 106 446
rect 0 100 1 101
rect 2 100 3 101
rect 3 100 4 101
rect 5 100 6 101
rect 0 101 6 105
rect 0 105 1 106
rect 2 105 3 106
rect 3 105 4 106
rect 5 105 6 106
rect 0 200 1 201
rect 2 200 3 201
rect 3 200 4 201
rect 5 200 6 201
rect 0 201 6 205
rect 0 205 1 206
rect 2 205 3 206
rect 3 205 4 206
rect 5 205 6 206
rect 260 300 261 301
rect 262 300 263 301
rect 263 300 264 301
rect 265 300 266 301
rect 260 301 266 305
rect 260 305 261 306
rect 262 305 263 306
rect 263 305 264 306
rect 265 305 266 306
rect 60 440 61 441
rect 62 440 63 441
rect 63 440 64 441
rect 65 440 66 441
rect 60 441 66 445
rect 60 445 61 446
rect 62 445 63 446
rect 63 445 64 446
rect 65 445 66 446
rect 340 0 341 1
rect 342 0 343 1
rect 343 0 344 1
rect 345 0 346 1
rect 340 1 346 5
rect 340 5 341 6
rect 342 5 343 6
rect 343 5 344 6
rect 345 5 346 6
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect 140 40 141 41
rect 142 40 143 41
rect 143 40 144 41
rect 145 40 146 41
rect 140 41 146 45
rect 140 45 141 46
rect 142 45 143 46
rect 143 45 144 46
rect 145 45 146 46
rect 520 260 521 261
rect 522 260 523 261
rect 523 260 524 261
rect 525 260 526 261
rect 520 261 526 265
rect 520 265 521 266
rect 522 265 523 266
rect 523 265 524 266
rect 525 265 526 266
rect 440 520 441 521
rect 442 520 443 521
rect 443 520 444 521
rect 445 520 446 521
rect 440 521 446 525
rect 440 525 441 526
rect 442 525 443 526
rect 443 525 444 526
rect 445 525 446 526
rect 160 460 161 461
rect 162 460 163 461
rect 163 460 164 461
rect 165 460 166 461
rect 160 461 166 465
rect 160 465 161 466
rect 162 465 163 466
rect 163 465 164 466
rect 165 465 166 466
rect 200 520 201 521
rect 202 520 203 521
rect 203 520 204 521
rect 205 520 206 521
rect 200 521 206 525
rect 200 525 201 526
rect 202 525 203 526
rect 203 525 204 526
rect 205 525 206 526
rect 540 300 541 301
rect 542 300 543 301
rect 543 300 544 301
rect 545 300 546 301
rect 540 301 546 305
rect 540 305 541 306
rect 542 305 543 306
rect 543 305 544 306
rect 545 305 546 306
rect 120 280 121 281
rect 122 280 123 281
rect 123 280 124 281
rect 125 280 126 281
rect 120 281 126 285
rect 120 285 121 286
rect 122 285 123 286
rect 123 285 124 286
rect 125 285 126 286
rect 100 320 101 321
rect 102 320 103 321
rect 103 320 104 321
rect 105 320 106 321
rect 100 321 106 325
rect 100 325 101 326
rect 102 325 103 326
rect 103 325 104 326
rect 105 325 106 326
rect 420 360 421 361
rect 422 360 423 361
rect 423 360 424 361
rect 425 360 426 361
rect 420 361 426 365
rect 420 365 421 366
rect 422 365 423 366
rect 423 365 424 366
rect 425 365 426 366
rect 360 100 361 101
rect 362 100 363 101
rect 363 100 364 101
rect 365 100 366 101
rect 360 101 366 105
rect 360 105 361 106
rect 362 105 363 106
rect 363 105 364 106
rect 365 105 366 106
rect 360 340 361 341
rect 362 340 363 341
rect 363 340 364 341
rect 365 340 366 341
rect 360 341 366 345
rect 360 345 361 346
rect 362 345 363 346
rect 363 345 364 346
rect 365 345 366 346
rect 320 240 321 241
rect 322 240 323 241
rect 323 240 324 241
rect 325 240 326 241
rect 320 241 326 245
rect 320 245 321 246
rect 322 245 323 246
rect 323 245 324 246
rect 325 245 326 246
rect 520 240 521 241
rect 522 240 523 241
rect 523 240 524 241
rect 525 240 526 241
rect 520 241 526 245
rect 520 245 521 246
rect 522 245 523 246
rect 523 245 524 246
rect 525 245 526 246
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect 280 480 281 481
rect 282 480 283 481
rect 283 480 284 481
rect 285 480 286 481
rect 280 481 286 485
rect 280 485 281 486
rect 282 485 283 486
rect 283 485 284 486
rect 285 485 286 486
rect 600 280 601 281
rect 602 280 603 281
rect 603 280 604 281
rect 605 280 606 281
rect 600 281 606 285
rect 600 285 601 286
rect 602 285 603 286
rect 603 285 604 286
rect 605 285 606 286
rect 300 360 301 361
rect 302 360 303 361
rect 303 360 304 361
rect 305 360 306 361
rect 300 361 306 365
rect 300 365 301 366
rect 302 365 303 366
rect 303 365 304 366
rect 305 365 306 366
rect 220 140 221 141
rect 222 140 223 141
rect 223 140 224 141
rect 225 140 226 141
rect 220 141 226 145
rect 220 145 221 146
rect 222 145 223 146
rect 223 145 224 146
rect 225 145 226 146
rect 200 100 201 101
rect 202 100 203 101
rect 203 100 204 101
rect 205 100 206 101
rect 200 101 206 105
rect 200 105 201 106
rect 202 105 203 106
rect 203 105 204 106
rect 205 105 206 106
rect 160 120 161 121
rect 162 120 163 121
rect 163 120 164 121
rect 165 120 166 121
rect 160 121 166 125
rect 160 125 161 126
rect 162 125 163 126
rect 163 125 164 126
rect 165 125 166 126
rect 440 380 441 381
rect 442 380 443 381
rect 443 380 444 381
rect 445 380 446 381
rect 440 381 446 385
rect 440 385 441 386
rect 442 385 443 386
rect 443 385 444 386
rect 445 385 446 386
rect 120 300 121 301
rect 122 300 123 301
rect 123 300 124 301
rect 125 300 126 301
rect 120 301 126 305
rect 120 305 121 306
rect 122 305 123 306
rect 123 305 124 306
rect 125 305 126 306
rect 220 360 221 361
rect 222 360 223 361
rect 223 360 224 361
rect 225 360 226 361
rect 220 361 226 365
rect 220 365 221 366
rect 222 365 223 366
rect 223 365 224 366
rect 225 365 226 366
rect 500 580 501 581
rect 502 580 503 581
rect 503 580 504 581
rect 505 580 506 581
rect 500 581 506 585
rect 500 585 501 586
rect 502 585 503 586
rect 503 585 504 586
rect 505 585 506 586
rect 500 220 501 221
rect 502 220 503 221
rect 503 220 504 221
rect 505 220 506 221
rect 500 221 506 225
rect 500 225 501 226
rect 502 225 503 226
rect 503 225 504 226
rect 505 225 506 226
rect 560 100 561 101
rect 562 100 563 101
rect 563 100 564 101
rect 565 100 566 101
rect 560 101 566 105
rect 560 105 561 106
rect 562 105 563 106
rect 563 105 564 106
rect 565 105 566 106
rect 180 440 181 441
rect 182 440 183 441
rect 183 440 184 441
rect 185 440 186 441
rect 180 441 186 445
rect 180 445 181 446
rect 182 445 183 446
rect 183 445 184 446
rect 185 445 186 446
rect 0 380 1 381
rect 2 380 3 381
rect 3 380 4 381
rect 5 380 6 381
rect 0 381 6 385
rect 0 385 1 386
rect 2 385 3 386
rect 3 385 4 386
rect 5 385 6 386
rect 200 20 201 21
rect 202 20 203 21
rect 203 20 204 21
rect 205 20 206 21
rect 200 21 206 25
rect 200 25 201 26
rect 202 25 203 26
rect 203 25 204 26
rect 205 25 206 26
rect 400 160 401 161
rect 402 160 403 161
rect 403 160 404 161
rect 405 160 406 161
rect 400 161 406 165
rect 400 165 401 166
rect 402 165 403 166
rect 403 165 404 166
rect 405 165 406 166
rect 460 220 461 221
rect 462 220 463 221
rect 463 220 464 221
rect 465 220 466 221
rect 460 221 466 225
rect 460 225 461 226
rect 462 225 463 226
rect 463 225 464 226
rect 465 225 466 226
rect 260 80 261 81
rect 262 80 263 81
rect 263 80 264 81
rect 265 80 266 81
rect 260 81 266 85
rect 260 85 261 86
rect 262 85 263 86
rect 263 85 264 86
rect 265 85 266 86
rect 180 620 181 621
rect 182 620 183 621
rect 183 620 184 621
rect 185 620 186 621
rect 180 621 186 625
rect 180 625 181 626
rect 182 625 183 626
rect 183 625 184 626
rect 185 625 186 626
rect 360 580 361 581
rect 362 580 363 581
rect 363 580 364 581
rect 365 580 366 581
rect 360 581 366 585
rect 360 585 361 586
rect 362 585 363 586
rect 363 585 364 586
rect 365 585 366 586
rect 480 60 481 61
rect 482 60 483 61
rect 483 60 484 61
rect 485 60 486 61
rect 480 61 486 65
rect 480 65 481 66
rect 482 65 483 66
rect 483 65 484 66
rect 485 65 486 66
rect 420 140 421 141
rect 422 140 423 141
rect 423 140 424 141
rect 425 140 426 141
rect 420 141 426 145
rect 420 145 421 146
rect 422 145 423 146
rect 423 145 424 146
rect 425 145 426 146
rect 560 300 561 301
rect 562 300 563 301
rect 563 300 564 301
rect 565 300 566 301
rect 560 301 566 305
rect 560 305 561 306
rect 562 305 563 306
rect 563 305 564 306
rect 565 305 566 306
rect 340 660 341 661
rect 342 660 343 661
rect 343 660 344 661
rect 345 660 346 661
rect 340 661 346 665
rect 340 665 341 666
rect 342 665 343 666
rect 343 665 344 666
rect 345 665 346 666
rect 200 140 201 141
rect 202 140 203 141
rect 203 140 204 141
rect 205 140 206 141
rect 200 141 206 145
rect 200 145 201 146
rect 202 145 203 146
rect 203 145 204 146
rect 205 145 206 146
rect 560 380 561 381
rect 562 380 563 381
rect 563 380 564 381
rect 565 380 566 381
rect 560 381 566 385
rect 560 385 561 386
rect 562 385 563 386
rect 563 385 564 386
rect 565 385 566 386
rect 40 380 41 381
rect 42 380 43 381
rect 43 380 44 381
rect 45 380 46 381
rect 40 381 46 385
rect 40 385 41 386
rect 42 385 43 386
rect 43 385 44 386
rect 45 385 46 386
rect 440 20 441 21
rect 442 20 443 21
rect 443 20 444 21
rect 445 20 446 21
rect 440 21 446 25
rect 440 25 441 26
rect 442 25 443 26
rect 443 25 444 26
rect 445 25 446 26
rect 600 220 601 221
rect 602 220 603 221
rect 603 220 604 221
rect 605 220 606 221
rect 600 221 606 225
rect 600 225 601 226
rect 602 225 603 226
rect 603 225 604 226
rect 605 225 606 226
rect 640 280 641 281
rect 642 280 643 281
rect 643 280 644 281
rect 645 280 646 281
rect 640 281 646 285
rect 640 285 641 286
rect 642 285 643 286
rect 643 285 644 286
rect 645 285 646 286
rect 520 380 521 381
rect 522 380 523 381
rect 523 380 524 381
rect 525 380 526 381
rect 520 381 526 385
rect 520 385 521 386
rect 522 385 523 386
rect 523 385 524 386
rect 525 385 526 386
rect 200 300 201 301
rect 202 300 203 301
rect 203 300 204 301
rect 205 300 206 301
rect 200 301 206 305
rect 200 305 201 306
rect 202 305 203 306
rect 203 305 204 306
rect 205 305 206 306
rect 440 300 441 301
rect 442 300 443 301
rect 443 300 444 301
rect 445 300 446 301
rect 440 301 446 305
rect 440 305 441 306
rect 442 305 443 306
rect 443 305 444 306
rect 445 305 446 306
rect 160 100 161 101
rect 162 100 163 101
rect 163 100 164 101
rect 165 100 166 101
rect 160 101 166 105
rect 160 105 161 106
rect 162 105 163 106
rect 163 105 164 106
rect 165 105 166 106
rect 100 140 101 141
rect 102 140 103 141
rect 103 140 104 141
rect 105 140 106 141
rect 100 141 106 145
rect 100 145 101 146
rect 102 145 103 146
rect 103 145 104 146
rect 105 145 106 146
rect 520 340 521 341
rect 522 340 523 341
rect 523 340 524 341
rect 525 340 526 341
rect 520 341 526 345
rect 520 345 521 346
rect 522 345 523 346
rect 523 345 524 346
rect 525 345 526 346
rect 220 0 221 1
rect 222 0 223 1
rect 223 0 224 1
rect 225 0 226 1
rect 220 1 226 5
rect 220 5 221 6
rect 222 5 223 6
rect 223 5 224 6
rect 225 5 226 6
rect 360 40 361 41
rect 362 40 363 41
rect 363 40 364 41
rect 365 40 366 41
rect 360 41 366 45
rect 360 45 361 46
rect 362 45 363 46
rect 363 45 364 46
rect 365 45 366 46
rect 20 320 21 321
rect 22 320 23 321
rect 23 320 24 321
rect 25 320 26 321
rect 20 321 26 325
rect 20 325 21 326
rect 22 325 23 326
rect 23 325 24 326
rect 25 325 26 326
rect 40 220 41 221
rect 42 220 43 221
rect 43 220 44 221
rect 45 220 46 221
rect 40 221 46 225
rect 40 225 41 226
rect 42 225 43 226
rect 43 225 44 226
rect 45 225 46 226
rect 440 580 441 581
rect 442 580 443 581
rect 443 580 444 581
rect 445 580 446 581
rect 440 581 446 585
rect 440 585 441 586
rect 442 585 443 586
rect 443 585 444 586
rect 445 585 446 586
rect 360 140 361 141
rect 362 140 363 141
rect 363 140 364 141
rect 365 140 366 141
rect 360 141 366 145
rect 360 145 361 146
rect 362 145 363 146
rect 363 145 364 146
rect 365 145 366 146
rect 400 640 401 641
rect 402 640 403 641
rect 403 640 404 641
rect 405 640 406 641
rect 400 641 406 645
rect 400 645 401 646
rect 402 645 403 646
rect 403 645 404 646
rect 405 645 406 646
rect 520 560 521 561
rect 522 560 523 561
rect 523 560 524 561
rect 525 560 526 561
rect 520 561 526 565
rect 520 565 521 566
rect 522 565 523 566
rect 523 565 524 566
rect 525 565 526 566
rect 20 340 21 341
rect 22 340 23 341
rect 23 340 24 341
rect 25 340 26 341
rect 20 341 26 345
rect 20 345 21 346
rect 22 345 23 346
rect 23 345 24 346
rect 25 345 26 346
rect 540 440 541 441
rect 542 440 543 441
rect 543 440 544 441
rect 545 440 546 441
rect 540 441 546 445
rect 540 445 541 446
rect 542 445 543 446
rect 543 445 544 446
rect 545 445 546 446
rect 420 320 421 321
rect 422 320 423 321
rect 423 320 424 321
rect 425 320 426 321
rect 420 321 426 325
rect 420 325 421 326
rect 422 325 423 326
rect 423 325 424 326
rect 425 325 426 326
rect 240 80 241 81
rect 242 80 243 81
rect 243 80 244 81
rect 245 80 246 81
rect 240 81 246 85
rect 240 85 241 86
rect 242 85 243 86
rect 243 85 244 86
rect 245 85 246 86
rect 560 520 561 521
rect 562 520 563 521
rect 563 520 564 521
rect 565 520 566 521
rect 560 521 566 525
rect 560 525 561 526
rect 562 525 563 526
rect 563 525 564 526
rect 565 525 566 526
rect 500 160 501 161
rect 502 160 503 161
rect 503 160 504 161
rect 505 160 506 161
rect 500 161 506 165
rect 500 165 501 166
rect 502 165 503 166
rect 503 165 504 166
rect 505 165 506 166
rect 80 420 81 421
rect 82 420 83 421
rect 83 420 84 421
rect 85 420 86 421
rect 80 421 86 425
rect 80 425 81 426
rect 82 425 83 426
rect 83 425 84 426
rect 85 425 86 426
rect 200 440 201 441
rect 202 440 203 441
rect 203 440 204 441
rect 205 440 206 441
rect 200 441 206 445
rect 200 445 201 446
rect 202 445 203 446
rect 203 445 204 446
rect 205 445 206 446
rect 80 500 81 501
rect 82 500 83 501
rect 83 500 84 501
rect 85 500 86 501
rect 80 501 86 505
rect 80 505 81 506
rect 82 505 83 506
rect 83 505 84 506
rect 85 505 86 506
rect 80 540 81 541
rect 82 540 83 541
rect 83 540 84 541
rect 85 540 86 541
rect 80 541 86 545
rect 80 545 81 546
rect 82 545 83 546
rect 83 545 84 546
rect 85 545 86 546
rect 60 360 61 361
rect 62 360 63 361
rect 63 360 64 361
rect 65 360 66 361
rect 60 361 66 365
rect 60 365 61 366
rect 62 365 63 366
rect 63 365 64 366
rect 65 365 66 366
rect 220 620 221 621
rect 222 620 223 621
rect 223 620 224 621
rect 225 620 226 621
rect 220 621 226 625
rect 220 625 221 626
rect 222 625 223 626
rect 223 625 224 626
rect 225 625 226 626
rect 320 420 321 421
rect 322 420 323 421
rect 323 420 324 421
rect 325 420 326 421
rect 320 421 326 425
rect 320 425 321 426
rect 322 425 323 426
rect 323 425 324 426
rect 325 425 326 426
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect 160 560 161 561
rect 162 560 163 561
rect 163 560 164 561
rect 165 560 166 561
rect 160 561 166 565
rect 160 565 161 566
rect 162 565 163 566
rect 163 565 164 566
rect 165 565 166 566
rect 440 200 441 201
rect 442 200 443 201
rect 443 200 444 201
rect 445 200 446 201
rect 440 201 446 205
rect 440 205 441 206
rect 442 205 443 206
rect 443 205 444 206
rect 445 205 446 206
rect 540 320 541 321
rect 542 320 543 321
rect 543 320 544 321
rect 545 320 546 321
rect 540 321 546 325
rect 540 325 541 326
rect 542 325 543 326
rect 543 325 544 326
rect 545 325 546 326
rect 620 300 621 301
rect 622 300 623 301
rect 623 300 624 301
rect 625 300 626 301
rect 620 301 626 305
rect 620 305 621 306
rect 622 305 623 306
rect 623 305 624 306
rect 625 305 626 306
rect 360 540 361 541
rect 362 540 363 541
rect 363 540 364 541
rect 365 540 366 541
rect 360 541 366 545
rect 360 545 361 546
rect 362 545 363 546
rect 363 545 364 546
rect 365 545 366 546
rect 300 660 301 661
rect 302 660 303 661
rect 303 660 304 661
rect 305 660 306 661
rect 300 661 306 665
rect 300 665 301 666
rect 302 665 303 666
rect 303 665 304 666
rect 305 665 306 666
rect 440 160 441 161
rect 442 160 443 161
rect 443 160 444 161
rect 445 160 446 161
rect 440 161 446 165
rect 440 165 441 166
rect 442 165 443 166
rect 443 165 444 166
rect 445 165 446 166
rect 20 360 21 361
rect 22 360 23 361
rect 23 360 24 361
rect 25 360 26 361
rect 20 361 26 365
rect 20 365 21 366
rect 22 365 23 366
rect 23 365 24 366
rect 25 365 26 366
rect 220 220 221 221
rect 222 220 223 221
rect 223 220 224 221
rect 225 220 226 221
rect 220 221 226 225
rect 220 225 221 226
rect 222 225 223 226
rect 223 225 224 226
rect 225 225 226 226
rect 160 360 161 361
rect 162 360 163 361
rect 163 360 164 361
rect 165 360 166 361
rect 160 361 166 365
rect 160 365 161 366
rect 162 365 163 366
rect 163 365 164 366
rect 165 365 166 366
rect 580 560 581 561
rect 582 560 583 561
rect 583 560 584 561
rect 585 560 586 561
rect 580 561 586 565
rect 580 565 581 566
rect 582 565 583 566
rect 583 565 584 566
rect 585 565 586 566
rect 80 240 81 241
rect 82 240 83 241
rect 83 240 84 241
rect 85 240 86 241
rect 80 241 86 245
rect 80 245 81 246
rect 82 245 83 246
rect 83 245 84 246
rect 85 245 86 246
rect 200 460 201 461
rect 202 460 203 461
rect 203 460 204 461
rect 205 460 206 461
rect 200 461 206 465
rect 200 465 201 466
rect 202 465 203 466
rect 203 465 204 466
rect 205 465 206 466
rect 540 460 541 461
rect 542 460 543 461
rect 543 460 544 461
rect 545 460 546 461
rect 540 461 546 465
rect 540 465 541 466
rect 542 465 543 466
rect 543 465 544 466
rect 545 465 546 466
rect 120 520 121 521
rect 122 520 123 521
rect 123 520 124 521
rect 125 520 126 521
rect 120 521 126 525
rect 120 525 121 526
rect 122 525 123 526
rect 123 525 124 526
rect 125 525 126 526
rect 500 0 501 1
rect 502 0 503 1
rect 503 0 504 1
rect 505 0 506 1
rect 500 1 506 5
rect 500 5 501 6
rect 502 5 503 6
rect 503 5 504 6
rect 505 5 506 6
rect 380 380 381 381
rect 382 380 383 381
rect 383 380 384 381
rect 385 380 386 381
rect 380 381 386 385
rect 380 385 381 386
rect 382 385 383 386
rect 383 385 384 386
rect 385 385 386 386
rect 480 120 481 121
rect 482 120 483 121
rect 483 120 484 121
rect 485 120 486 121
rect 480 121 486 125
rect 480 125 481 126
rect 482 125 483 126
rect 483 125 484 126
rect 485 125 486 126
rect 300 260 301 261
rect 302 260 303 261
rect 303 260 304 261
rect 305 260 306 261
rect 300 261 306 265
rect 300 265 301 266
rect 302 265 303 266
rect 303 265 304 266
rect 305 265 306 266
rect 560 280 561 281
rect 562 280 563 281
rect 563 280 564 281
rect 565 280 566 281
rect 560 281 566 285
rect 560 285 561 286
rect 562 285 563 286
rect 563 285 564 286
rect 565 285 566 286
rect 340 580 341 581
rect 342 580 343 581
rect 343 580 344 581
rect 345 580 346 581
rect 340 581 346 585
rect 340 585 341 586
rect 342 585 343 586
rect 343 585 344 586
rect 345 585 346 586
rect 280 180 281 181
rect 282 180 283 181
rect 283 180 284 181
rect 285 180 286 181
rect 280 181 286 185
rect 280 185 281 186
rect 282 185 283 186
rect 283 185 284 186
rect 285 185 286 186
rect 480 220 481 221
rect 482 220 483 221
rect 483 220 484 221
rect 485 220 486 221
rect 480 221 486 225
rect 480 225 481 226
rect 482 225 483 226
rect 483 225 484 226
rect 485 225 486 226
rect 180 360 181 361
rect 182 360 183 361
rect 183 360 184 361
rect 185 360 186 361
rect 180 361 186 365
rect 180 365 181 366
rect 182 365 183 366
rect 183 365 184 366
rect 185 365 186 366
rect 80 200 81 201
rect 82 200 83 201
rect 83 200 84 201
rect 85 200 86 201
rect 80 201 86 205
rect 80 205 81 206
rect 82 205 83 206
rect 83 205 84 206
rect 85 205 86 206
rect 380 240 381 241
rect 382 240 383 241
rect 383 240 384 241
rect 385 240 386 241
rect 380 241 386 245
rect 380 245 381 246
rect 382 245 383 246
rect 383 245 384 246
rect 385 245 386 246
rect 0 360 1 361
rect 2 360 3 361
rect 3 360 4 361
rect 5 360 6 361
rect 0 361 6 365
rect 0 365 1 366
rect 2 365 3 366
rect 3 365 4 366
rect 5 365 6 366
rect 320 300 321 301
rect 322 300 323 301
rect 323 300 324 301
rect 325 300 326 301
rect 320 301 326 305
rect 320 305 321 306
rect 322 305 323 306
rect 323 305 324 306
rect 325 305 326 306
rect 420 520 421 521
rect 422 520 423 521
rect 423 520 424 521
rect 425 520 426 521
rect 420 521 426 525
rect 420 525 421 526
rect 422 525 423 526
rect 423 525 424 526
rect 425 525 426 526
rect 380 520 381 521
rect 382 520 383 521
rect 383 520 384 521
rect 385 520 386 521
rect 380 521 386 525
rect 380 525 381 526
rect 382 525 383 526
rect 383 525 384 526
rect 385 525 386 526
rect 40 200 41 201
rect 42 200 43 201
rect 43 200 44 201
rect 45 200 46 201
rect 40 201 46 205
rect 40 205 41 206
rect 42 205 43 206
rect 43 205 44 206
rect 45 205 46 206
rect 280 40 281 41
rect 282 40 283 41
rect 283 40 284 41
rect 285 40 286 41
rect 280 41 286 45
rect 280 45 281 46
rect 282 45 283 46
rect 283 45 284 46
rect 285 45 286 46
rect 280 640 281 641
rect 282 640 283 641
rect 283 640 284 641
rect 285 640 286 641
rect 280 641 286 645
rect 280 645 281 646
rect 282 645 283 646
rect 283 645 284 646
rect 285 645 286 646
rect 180 140 181 141
rect 182 140 183 141
rect 183 140 184 141
rect 185 140 186 141
rect 180 141 186 145
rect 180 145 181 146
rect 182 145 183 146
rect 183 145 184 146
rect 185 145 186 146
rect 280 280 281 281
rect 282 280 283 281
rect 283 280 284 281
rect 285 280 286 281
rect 280 281 286 285
rect 280 285 281 286
rect 282 285 283 286
rect 283 285 284 286
rect 285 285 286 286
rect 320 580 321 581
rect 322 580 323 581
rect 323 580 324 581
rect 325 580 326 581
rect 320 581 326 585
rect 320 585 321 586
rect 322 585 323 586
rect 323 585 324 586
rect 325 585 326 586
rect 140 480 141 481
rect 142 480 143 481
rect 143 480 144 481
rect 145 480 146 481
rect 140 481 146 485
rect 140 485 141 486
rect 142 485 143 486
rect 143 485 144 486
rect 145 485 146 486
rect 140 460 141 461
rect 142 460 143 461
rect 143 460 144 461
rect 145 460 146 461
rect 140 461 146 465
rect 140 465 141 466
rect 142 465 143 466
rect 143 465 144 466
rect 145 465 146 466
rect 60 340 61 341
rect 62 340 63 341
rect 63 340 64 341
rect 65 340 66 341
rect 60 341 66 345
rect 60 345 61 346
rect 62 345 63 346
rect 63 345 64 346
rect 65 345 66 346
rect 100 180 101 181
rect 102 180 103 181
rect 103 180 104 181
rect 105 180 106 181
rect 100 181 106 185
rect 100 185 101 186
rect 102 185 103 186
rect 103 185 104 186
rect 105 185 106 186
rect 620 480 621 481
rect 622 480 623 481
rect 623 480 624 481
rect 625 480 626 481
rect 620 481 626 485
rect 620 485 621 486
rect 622 485 623 486
rect 623 485 624 486
rect 625 485 626 486
rect 400 180 401 181
rect 402 180 403 181
rect 403 180 404 181
rect 405 180 406 181
rect 400 181 406 185
rect 400 185 401 186
rect 402 185 403 186
rect 403 185 404 186
rect 405 185 406 186
rect 240 640 241 641
rect 242 640 243 641
rect 243 640 244 641
rect 245 640 246 641
rect 240 641 246 645
rect 240 645 241 646
rect 242 645 243 646
rect 243 645 244 646
rect 245 645 246 646
rect 300 240 301 241
rect 302 240 303 241
rect 303 240 304 241
rect 305 240 306 241
rect 300 241 306 245
rect 300 245 301 246
rect 302 245 303 246
rect 303 245 304 246
rect 305 245 306 246
rect 320 200 321 201
rect 322 200 323 201
rect 323 200 324 201
rect 325 200 326 201
rect 320 201 326 205
rect 320 205 321 206
rect 322 205 323 206
rect 323 205 324 206
rect 325 205 326 206
rect 80 100 81 101
rect 82 100 83 101
rect 83 100 84 101
rect 85 100 86 101
rect 80 101 86 105
rect 80 105 81 106
rect 82 105 83 106
rect 83 105 84 106
rect 85 105 86 106
rect 380 200 381 201
rect 382 200 383 201
rect 383 200 384 201
rect 385 200 386 201
rect 380 201 386 205
rect 380 205 381 206
rect 382 205 383 206
rect 383 205 384 206
rect 385 205 386 206
rect 500 40 501 41
rect 502 40 503 41
rect 503 40 504 41
rect 505 40 506 41
rect 500 41 506 45
rect 500 45 501 46
rect 502 45 503 46
rect 503 45 504 46
rect 505 45 506 46
rect 340 60 341 61
rect 342 60 343 61
rect 343 60 344 61
rect 345 60 346 61
rect 340 61 346 65
rect 340 65 341 66
rect 342 65 343 66
rect 343 65 344 66
rect 345 65 346 66
rect 360 360 361 361
rect 362 360 363 361
rect 363 360 364 361
rect 365 360 366 361
rect 360 361 366 365
rect 360 365 361 366
rect 362 365 363 366
rect 363 365 364 366
rect 365 365 366 366
rect 580 400 581 401
rect 582 400 583 401
rect 583 400 584 401
rect 585 400 586 401
rect 580 401 586 405
rect 580 405 581 406
rect 582 405 583 406
rect 583 405 584 406
rect 585 405 586 406
rect 200 380 201 381
rect 202 380 203 381
rect 203 380 204 381
rect 205 380 206 381
rect 200 381 206 385
rect 200 385 201 386
rect 202 385 203 386
rect 203 385 204 386
rect 205 385 206 386
rect 120 600 121 601
rect 122 600 123 601
rect 123 600 124 601
rect 125 600 126 601
rect 120 601 126 605
rect 120 605 121 606
rect 122 605 123 606
rect 123 605 124 606
rect 125 605 126 606
rect 40 320 41 321
rect 42 320 43 321
rect 43 320 44 321
rect 45 320 46 321
rect 40 321 46 325
rect 40 325 41 326
rect 42 325 43 326
rect 43 325 44 326
rect 45 325 46 326
rect 60 180 61 181
rect 62 180 63 181
rect 63 180 64 181
rect 65 180 66 181
rect 60 181 66 185
rect 60 185 61 186
rect 62 185 63 186
rect 63 185 64 186
rect 65 185 66 186
rect 320 600 321 601
rect 322 600 323 601
rect 323 600 324 601
rect 325 600 326 601
rect 320 601 326 605
rect 320 605 321 606
rect 322 605 323 606
rect 323 605 324 606
rect 325 605 326 606
rect 100 80 101 81
rect 102 80 103 81
rect 103 80 104 81
rect 105 80 106 81
rect 100 81 106 85
rect 100 85 101 86
rect 102 85 103 86
rect 103 85 104 86
rect 105 85 106 86
rect 180 180 181 181
rect 182 180 183 181
rect 183 180 184 181
rect 185 180 186 181
rect 180 181 186 185
rect 180 185 181 186
rect 182 185 183 186
rect 183 185 184 186
rect 185 185 186 186
rect 200 420 201 421
rect 202 420 203 421
rect 203 420 204 421
rect 205 420 206 421
rect 200 421 206 425
rect 200 425 201 426
rect 202 425 203 426
rect 203 425 204 426
rect 205 425 206 426
rect 420 100 421 101
rect 422 100 423 101
rect 423 100 424 101
rect 425 100 426 101
rect 420 101 426 105
rect 420 105 421 106
rect 422 105 423 106
rect 423 105 424 106
rect 425 105 426 106
rect 500 540 501 541
rect 502 540 503 541
rect 503 540 504 541
rect 505 540 506 541
rect 500 541 506 545
rect 500 545 501 546
rect 502 545 503 546
rect 503 545 504 546
rect 505 545 506 546
rect 580 420 581 421
rect 582 420 583 421
rect 583 420 584 421
rect 585 420 586 421
rect 580 421 586 425
rect 580 425 581 426
rect 582 425 583 426
rect 583 425 584 426
rect 585 425 586 426
rect 560 200 561 201
rect 562 200 563 201
rect 563 200 564 201
rect 565 200 566 201
rect 560 201 566 205
rect 560 205 561 206
rect 562 205 563 206
rect 563 205 564 206
rect 565 205 566 206
rect 540 420 541 421
rect 542 420 543 421
rect 543 420 544 421
rect 545 420 546 421
rect 540 421 546 425
rect 540 425 541 426
rect 542 425 543 426
rect 543 425 544 426
rect 545 425 546 426
rect 300 320 301 321
rect 302 320 303 321
rect 303 320 304 321
rect 305 320 306 321
rect 300 321 306 325
rect 300 325 301 326
rect 302 325 303 326
rect 303 325 304 326
rect 305 325 306 326
rect 260 400 261 401
rect 262 400 263 401
rect 263 400 264 401
rect 265 400 266 401
rect 260 401 266 405
rect 260 405 261 406
rect 262 405 263 406
rect 263 405 264 406
rect 265 405 266 406
rect 320 320 321 321
rect 322 320 323 321
rect 323 320 324 321
rect 325 320 326 321
rect 320 321 326 325
rect 320 325 321 326
rect 322 325 323 326
rect 323 325 324 326
rect 325 325 326 326
rect 220 540 221 541
rect 222 540 223 541
rect 223 540 224 541
rect 225 540 226 541
rect 220 541 226 545
rect 220 545 221 546
rect 222 545 223 546
rect 223 545 224 546
rect 225 545 226 546
rect 420 380 421 381
rect 422 380 423 381
rect 423 380 424 381
rect 425 380 426 381
rect 420 381 426 385
rect 420 385 421 386
rect 422 385 423 386
rect 423 385 424 386
rect 425 385 426 386
rect 300 80 301 81
rect 302 80 303 81
rect 303 80 304 81
rect 305 80 306 81
rect 300 81 306 85
rect 300 85 301 86
rect 302 85 303 86
rect 303 85 304 86
rect 305 85 306 86
rect 160 380 161 381
rect 162 380 163 381
rect 163 380 164 381
rect 165 380 166 381
rect 160 381 166 385
rect 160 385 161 386
rect 162 385 163 386
rect 163 385 164 386
rect 165 385 166 386
rect 160 500 161 501
rect 162 500 163 501
rect 163 500 164 501
rect 165 500 166 501
rect 160 501 166 505
rect 160 505 161 506
rect 162 505 163 506
rect 163 505 164 506
rect 165 505 166 506
rect 480 500 481 501
rect 482 500 483 501
rect 483 500 484 501
rect 485 500 486 501
rect 480 501 486 505
rect 480 505 481 506
rect 482 505 483 506
rect 483 505 484 506
rect 485 505 486 506
rect 60 80 61 81
rect 62 80 63 81
rect 63 80 64 81
rect 65 80 66 81
rect 60 81 66 85
rect 60 85 61 86
rect 62 85 63 86
rect 63 85 64 86
rect 65 85 66 86
rect 480 420 481 421
rect 482 420 483 421
rect 483 420 484 421
rect 485 420 486 421
rect 480 421 486 425
rect 480 425 481 426
rect 482 425 483 426
rect 483 425 484 426
rect 485 425 486 426
rect 380 400 381 401
rect 382 400 383 401
rect 383 400 384 401
rect 385 400 386 401
rect 380 401 386 405
rect 380 405 381 406
rect 382 405 383 406
rect 383 405 384 406
rect 385 405 386 406
rect 560 140 561 141
rect 562 140 563 141
rect 563 140 564 141
rect 565 140 566 141
rect 560 141 566 145
rect 560 145 561 146
rect 562 145 563 146
rect 563 145 564 146
rect 565 145 566 146
rect 200 540 201 541
rect 202 540 203 541
rect 203 540 204 541
rect 205 540 206 541
rect 200 541 206 545
rect 200 545 201 546
rect 202 545 203 546
rect 203 545 204 546
rect 205 545 206 546
rect 440 180 441 181
rect 442 180 443 181
rect 443 180 444 181
rect 445 180 446 181
rect 440 181 446 185
rect 440 185 441 186
rect 442 185 443 186
rect 443 185 444 186
rect 445 185 446 186
rect 620 420 621 421
rect 622 420 623 421
rect 623 420 624 421
rect 625 420 626 421
rect 620 421 626 425
rect 620 425 621 426
rect 622 425 623 426
rect 623 425 624 426
rect 625 425 626 426
rect 180 260 181 261
rect 182 260 183 261
rect 183 260 184 261
rect 185 260 186 261
rect 180 261 186 265
rect 180 265 181 266
rect 182 265 183 266
rect 183 265 184 266
rect 185 265 186 266
rect 220 660 221 661
rect 222 660 223 661
rect 223 660 224 661
rect 225 660 226 661
rect 220 661 226 665
rect 220 665 221 666
rect 222 665 223 666
rect 223 665 224 666
rect 225 665 226 666
rect 360 420 361 421
rect 362 420 363 421
rect 363 420 364 421
rect 365 420 366 421
rect 360 421 366 425
rect 360 425 361 426
rect 362 425 363 426
rect 363 425 364 426
rect 365 425 366 426
rect 120 60 121 61
rect 122 60 123 61
rect 123 60 124 61
rect 125 60 126 61
rect 120 61 126 65
rect 120 65 121 66
rect 122 65 123 66
rect 123 65 124 66
rect 125 65 126 66
rect 660 440 661 441
rect 662 440 663 441
rect 663 440 664 441
rect 665 440 666 441
rect 660 441 666 445
rect 660 445 661 446
rect 662 445 663 446
rect 663 445 664 446
rect 665 445 666 446
rect 200 340 201 341
rect 202 340 203 341
rect 203 340 204 341
rect 205 340 206 341
rect 200 341 206 345
rect 200 345 201 346
rect 202 345 203 346
rect 203 345 204 346
rect 205 345 206 346
rect 540 40 541 41
rect 542 40 543 41
rect 543 40 544 41
rect 545 40 546 41
rect 540 41 546 45
rect 540 45 541 46
rect 542 45 543 46
rect 543 45 544 46
rect 545 45 546 46
rect 520 0 521 1
rect 522 0 523 1
rect 523 0 524 1
rect 525 0 526 1
rect 520 1 526 5
rect 520 5 521 6
rect 522 5 523 6
rect 523 5 524 6
rect 525 5 526 6
rect 580 460 581 461
rect 582 460 583 461
rect 583 460 584 461
rect 585 460 586 461
rect 580 461 586 465
rect 580 465 581 466
rect 582 465 583 466
rect 583 465 584 466
rect 585 465 586 466
rect 180 160 181 161
rect 182 160 183 161
rect 183 160 184 161
rect 185 160 186 161
rect 180 161 186 165
rect 180 165 181 166
rect 182 165 183 166
rect 183 165 184 166
rect 185 165 186 166
rect 540 120 541 121
rect 542 120 543 121
rect 543 120 544 121
rect 545 120 546 121
rect 540 121 546 125
rect 540 125 541 126
rect 542 125 543 126
rect 543 125 544 126
rect 545 125 546 126
rect 420 40 421 41
rect 422 40 423 41
rect 423 40 424 41
rect 425 40 426 41
rect 420 41 426 45
rect 420 45 421 46
rect 422 45 423 46
rect 423 45 424 46
rect 425 45 426 46
rect 400 440 401 441
rect 402 440 403 441
rect 403 440 404 441
rect 405 440 406 441
rect 400 441 406 445
rect 400 445 401 446
rect 402 445 403 446
rect 403 445 404 446
rect 405 445 406 446
rect 140 360 141 361
rect 142 360 143 361
rect 143 360 144 361
rect 145 360 146 361
rect 140 361 146 365
rect 140 365 141 366
rect 142 365 143 366
rect 143 365 144 366
rect 145 365 146 366
rect 440 240 441 241
rect 442 240 443 241
rect 443 240 444 241
rect 445 240 446 241
rect 440 241 446 245
rect 440 245 441 246
rect 442 245 443 246
rect 443 245 444 246
rect 445 245 446 246
rect 360 200 361 201
rect 362 200 363 201
rect 363 200 364 201
rect 365 200 366 201
rect 360 201 366 205
rect 360 205 361 206
rect 362 205 363 206
rect 363 205 364 206
rect 365 205 366 206
rect 440 560 441 561
rect 442 560 443 561
rect 443 560 444 561
rect 445 560 446 561
rect 440 561 446 565
rect 440 565 441 566
rect 442 565 443 566
rect 443 565 444 566
rect 445 565 446 566
rect 180 280 181 281
rect 182 280 183 281
rect 183 280 184 281
rect 185 280 186 281
rect 180 281 186 285
rect 180 285 181 286
rect 182 285 183 286
rect 183 285 184 286
rect 185 285 186 286
rect 540 160 541 161
rect 542 160 543 161
rect 543 160 544 161
rect 545 160 546 161
rect 540 161 546 165
rect 540 165 541 166
rect 542 165 543 166
rect 543 165 544 166
rect 545 165 546 166
rect 80 360 81 361
rect 82 360 83 361
rect 83 360 84 361
rect 85 360 86 361
rect 80 361 86 365
rect 80 365 81 366
rect 82 365 83 366
rect 83 365 84 366
rect 85 365 86 366
rect 240 340 241 341
rect 242 340 243 341
rect 243 340 244 341
rect 245 340 246 341
rect 240 341 246 345
rect 240 345 241 346
rect 242 345 243 346
rect 243 345 244 346
rect 245 345 246 346
rect 140 340 141 341
rect 142 340 143 341
rect 143 340 144 341
rect 145 340 146 341
rect 140 341 146 345
rect 140 345 141 346
rect 142 345 143 346
rect 143 345 144 346
rect 145 345 146 346
rect 240 560 241 561
rect 242 560 243 561
rect 243 560 244 561
rect 245 560 246 561
rect 240 561 246 565
rect 240 565 241 566
rect 242 565 243 566
rect 243 565 244 566
rect 245 565 246 566
rect 300 40 301 41
rect 302 40 303 41
rect 303 40 304 41
rect 305 40 306 41
rect 300 41 306 45
rect 300 45 301 46
rect 302 45 303 46
rect 303 45 304 46
rect 305 45 306 46
rect 180 200 181 201
rect 182 200 183 201
rect 183 200 184 201
rect 185 200 186 201
rect 180 201 186 205
rect 180 205 181 206
rect 182 205 183 206
rect 183 205 184 206
rect 185 205 186 206
rect 260 460 261 461
rect 262 460 263 461
rect 263 460 264 461
rect 265 460 266 461
rect 260 461 266 465
rect 260 465 261 466
rect 262 465 263 466
rect 263 465 264 466
rect 265 465 266 466
rect 420 120 421 121
rect 422 120 423 121
rect 423 120 424 121
rect 425 120 426 121
rect 420 121 426 125
rect 420 125 421 126
rect 422 125 423 126
rect 423 125 424 126
rect 425 125 426 126
rect 540 0 541 1
rect 542 0 543 1
rect 543 0 544 1
rect 545 0 546 1
rect 540 1 546 5
rect 540 5 541 6
rect 542 5 543 6
rect 543 5 544 6
rect 545 5 546 6
rect 280 100 281 101
rect 282 100 283 101
rect 283 100 284 101
rect 285 100 286 101
rect 280 101 286 105
rect 280 105 281 106
rect 282 105 283 106
rect 283 105 284 106
rect 285 105 286 106
rect 140 200 141 201
rect 142 200 143 201
rect 143 200 144 201
rect 145 200 146 201
rect 140 201 146 205
rect 140 205 141 206
rect 142 205 143 206
rect 143 205 144 206
rect 145 205 146 206
rect 380 0 381 1
rect 382 0 383 1
rect 383 0 384 1
rect 385 0 386 1
rect 380 1 386 5
rect 380 5 381 6
rect 382 5 383 6
rect 383 5 384 6
rect 385 5 386 6
rect 540 400 541 401
rect 542 400 543 401
rect 543 400 544 401
rect 545 400 546 401
rect 540 401 546 405
rect 540 405 541 406
rect 542 405 543 406
rect 543 405 544 406
rect 545 405 546 406
rect 460 40 461 41
rect 462 40 463 41
rect 463 40 464 41
rect 465 40 466 41
rect 460 41 466 45
rect 460 45 461 46
rect 462 45 463 46
rect 463 45 464 46
rect 465 45 466 46
rect 380 340 381 341
rect 382 340 383 341
rect 383 340 384 341
rect 385 340 386 341
rect 380 341 386 345
rect 380 345 381 346
rect 382 345 383 346
rect 383 345 384 346
rect 385 345 386 346
rect 520 440 521 441
rect 522 440 523 441
rect 523 440 524 441
rect 525 440 526 441
rect 520 441 526 445
rect 520 445 521 446
rect 522 445 523 446
rect 523 445 524 446
rect 525 445 526 446
rect 300 100 301 101
rect 302 100 303 101
rect 303 100 304 101
rect 305 100 306 101
rect 300 101 306 105
rect 300 105 301 106
rect 302 105 303 106
rect 303 105 304 106
rect 305 105 306 106
rect 240 200 241 201
rect 242 200 243 201
rect 243 200 244 201
rect 245 200 246 201
rect 240 201 246 205
rect 240 205 241 206
rect 242 205 243 206
rect 243 205 244 206
rect 245 205 246 206
rect 500 20 501 21
rect 502 20 503 21
rect 503 20 504 21
rect 505 20 506 21
rect 500 21 506 25
rect 500 25 501 26
rect 502 25 503 26
rect 503 25 504 26
rect 505 25 506 26
rect 60 540 61 541
rect 62 540 63 541
rect 63 540 64 541
rect 65 540 66 541
rect 60 541 66 545
rect 60 545 61 546
rect 62 545 63 546
rect 63 545 64 546
rect 65 545 66 546
rect 160 280 161 281
rect 162 280 163 281
rect 163 280 164 281
rect 165 280 166 281
rect 160 281 166 285
rect 160 285 161 286
rect 162 285 163 286
rect 163 285 164 286
rect 165 285 166 286
rect 400 560 401 561
rect 402 560 403 561
rect 403 560 404 561
rect 405 560 406 561
rect 400 561 406 565
rect 400 565 401 566
rect 402 565 403 566
rect 403 565 404 566
rect 405 565 406 566
rect 500 320 501 321
rect 502 320 503 321
rect 503 320 504 321
rect 505 320 506 321
rect 500 321 506 325
rect 500 325 501 326
rect 502 325 503 326
rect 503 325 504 326
rect 505 325 506 326
rect 120 480 121 481
rect 122 480 123 481
rect 123 480 124 481
rect 125 480 126 481
rect 120 481 126 485
rect 120 485 121 486
rect 122 485 123 486
rect 123 485 124 486
rect 125 485 126 486
rect 120 580 121 581
rect 122 580 123 581
rect 123 580 124 581
rect 125 580 126 581
rect 120 581 126 585
rect 120 585 121 586
rect 122 585 123 586
rect 123 585 124 586
rect 125 585 126 586
rect 520 600 521 601
rect 522 600 523 601
rect 523 600 524 601
rect 525 600 526 601
rect 520 601 526 605
rect 520 605 521 606
rect 522 605 523 606
rect 523 605 524 606
rect 525 605 526 606
rect 540 520 541 521
rect 542 520 543 521
rect 543 520 544 521
rect 545 520 546 521
rect 540 521 546 525
rect 540 525 541 526
rect 542 525 543 526
rect 543 525 544 526
rect 545 525 546 526
rect 320 40 321 41
rect 322 40 323 41
rect 323 40 324 41
rect 325 40 326 41
rect 320 41 326 45
rect 320 45 321 46
rect 322 45 323 46
rect 323 45 324 46
rect 325 45 326 46
rect 360 560 361 561
rect 362 560 363 561
rect 363 560 364 561
rect 365 560 366 561
rect 360 561 366 565
rect 360 565 361 566
rect 362 565 363 566
rect 363 565 364 566
rect 365 565 366 566
rect 300 580 301 581
rect 302 580 303 581
rect 303 580 304 581
rect 305 580 306 581
rect 300 581 306 585
rect 300 585 301 586
rect 302 585 303 586
rect 303 585 304 586
rect 305 585 306 586
rect 440 360 441 361
rect 442 360 443 361
rect 443 360 444 361
rect 445 360 446 361
rect 440 361 446 365
rect 440 365 441 366
rect 442 365 443 366
rect 443 365 444 366
rect 445 365 446 366
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect 420 300 421 301
rect 422 300 423 301
rect 423 300 424 301
rect 425 300 426 301
rect 420 301 426 305
rect 420 305 421 306
rect 422 305 423 306
rect 423 305 424 306
rect 425 305 426 306
rect 360 600 361 601
rect 362 600 363 601
rect 363 600 364 601
rect 365 600 366 601
rect 360 601 366 605
rect 360 605 361 606
rect 362 605 363 606
rect 363 605 364 606
rect 365 605 366 606
rect 440 260 441 261
rect 442 260 443 261
rect 443 260 444 261
rect 445 260 446 261
rect 440 261 446 265
rect 440 265 441 266
rect 442 265 443 266
rect 443 265 444 266
rect 445 265 446 266
rect 300 160 301 161
rect 302 160 303 161
rect 303 160 304 161
rect 305 160 306 161
rect 300 161 306 165
rect 300 165 301 166
rect 302 165 303 166
rect 303 165 304 166
rect 305 165 306 166
rect 220 300 221 301
rect 222 300 223 301
rect 223 300 224 301
rect 225 300 226 301
rect 220 301 226 305
rect 220 305 221 306
rect 222 305 223 306
rect 223 305 224 306
rect 225 305 226 306
rect 440 80 441 81
rect 442 80 443 81
rect 443 80 444 81
rect 445 80 446 81
rect 440 81 446 85
rect 440 85 441 86
rect 442 85 443 86
rect 443 85 444 86
rect 445 85 446 86
rect 460 620 461 621
rect 462 620 463 621
rect 463 620 464 621
rect 465 620 466 621
rect 460 621 466 625
rect 460 625 461 626
rect 462 625 463 626
rect 463 625 464 626
rect 465 625 466 626
rect 200 180 201 181
rect 202 180 203 181
rect 203 180 204 181
rect 205 180 206 181
rect 200 181 206 185
rect 200 185 201 186
rect 202 185 203 186
rect 203 185 204 186
rect 205 185 206 186
rect 40 500 41 501
rect 42 500 43 501
rect 43 500 44 501
rect 45 500 46 501
rect 40 501 46 505
rect 40 505 41 506
rect 42 505 43 506
rect 43 505 44 506
rect 45 505 46 506
rect 420 540 421 541
rect 422 540 423 541
rect 423 540 424 541
rect 425 540 426 541
rect 420 541 426 545
rect 420 545 421 546
rect 422 545 423 546
rect 423 545 424 546
rect 425 545 426 546
rect 140 580 141 581
rect 142 580 143 581
rect 143 580 144 581
rect 145 580 146 581
rect 140 581 146 585
rect 140 585 141 586
rect 142 585 143 586
rect 143 585 144 586
rect 145 585 146 586
rect 320 140 321 141
rect 322 140 323 141
rect 323 140 324 141
rect 325 140 326 141
rect 320 141 326 145
rect 320 145 321 146
rect 322 145 323 146
rect 323 145 324 146
rect 325 145 326 146
rect 220 200 221 201
rect 222 200 223 201
rect 223 200 224 201
rect 225 200 226 201
rect 220 201 226 205
rect 220 205 221 206
rect 222 205 223 206
rect 223 205 224 206
rect 225 205 226 206
rect 120 40 121 41
rect 122 40 123 41
rect 123 40 124 41
rect 125 40 126 41
rect 120 41 126 45
rect 120 45 121 46
rect 122 45 123 46
rect 123 45 124 46
rect 125 45 126 46
rect 60 140 61 141
rect 62 140 63 141
rect 63 140 64 141
rect 65 140 66 141
rect 60 141 66 145
rect 60 145 61 146
rect 62 145 63 146
rect 63 145 64 146
rect 65 145 66 146
rect 220 640 221 641
rect 222 640 223 641
rect 223 640 224 641
rect 225 640 226 641
rect 220 641 226 645
rect 220 645 221 646
rect 222 645 223 646
rect 223 645 224 646
rect 225 645 226 646
rect 600 480 601 481
rect 602 480 603 481
rect 603 480 604 481
rect 605 480 606 481
rect 600 481 606 485
rect 600 485 601 486
rect 602 485 603 486
rect 603 485 604 486
rect 605 485 606 486
rect 540 560 541 561
rect 542 560 543 561
rect 543 560 544 561
rect 545 560 546 561
rect 540 561 546 565
rect 540 565 541 566
rect 542 565 543 566
rect 543 565 544 566
rect 545 565 546 566
rect 280 220 281 221
rect 282 220 283 221
rect 283 220 284 221
rect 285 220 286 221
rect 280 221 286 225
rect 280 225 281 226
rect 282 225 283 226
rect 283 225 284 226
rect 285 225 286 226
rect 0 340 1 341
rect 2 340 3 341
rect 3 340 4 341
rect 5 340 6 341
rect 0 341 6 345
rect 0 345 1 346
rect 2 345 3 346
rect 3 345 4 346
rect 5 345 6 346
rect 440 420 441 421
rect 442 420 443 421
rect 443 420 444 421
rect 445 420 446 421
rect 440 421 446 425
rect 440 425 441 426
rect 442 425 443 426
rect 443 425 444 426
rect 445 425 446 426
rect 480 300 481 301
rect 482 300 483 301
rect 483 300 484 301
rect 485 300 486 301
rect 480 301 486 305
rect 480 305 481 306
rect 482 305 483 306
rect 483 305 484 306
rect 485 305 486 306
rect 0 480 1 481
rect 2 480 3 481
rect 3 480 4 481
rect 5 480 6 481
rect 0 481 6 485
rect 0 485 1 486
rect 2 485 3 486
rect 3 485 4 486
rect 5 485 6 486
rect 520 220 521 221
rect 522 220 523 221
rect 523 220 524 221
rect 525 220 526 221
rect 520 221 526 225
rect 520 225 521 226
rect 522 225 523 226
rect 523 225 524 226
rect 525 225 526 226
rect 260 20 261 21
rect 262 20 263 21
rect 263 20 264 21
rect 265 20 266 21
rect 260 21 266 25
rect 260 25 261 26
rect 262 25 263 26
rect 263 25 264 26
rect 265 25 266 26
rect 460 160 461 161
rect 462 160 463 161
rect 463 160 464 161
rect 465 160 466 161
rect 460 161 466 165
rect 460 165 461 166
rect 462 165 463 166
rect 463 165 464 166
rect 465 165 466 166
rect 360 80 361 81
rect 362 80 363 81
rect 363 80 364 81
rect 365 80 366 81
rect 360 81 366 85
rect 360 85 361 86
rect 362 85 363 86
rect 363 85 364 86
rect 365 85 366 86
rect 340 420 341 421
rect 342 420 343 421
rect 343 420 344 421
rect 345 420 346 421
rect 340 421 346 425
rect 340 425 341 426
rect 342 425 343 426
rect 343 425 344 426
rect 345 425 346 426
rect 300 120 301 121
rect 302 120 303 121
rect 303 120 304 121
rect 305 120 306 121
rect 300 121 306 125
rect 300 125 301 126
rect 302 125 303 126
rect 303 125 304 126
rect 305 125 306 126
rect 660 220 661 221
rect 662 220 663 221
rect 663 220 664 221
rect 665 220 666 221
rect 660 221 666 225
rect 660 225 661 226
rect 662 225 663 226
rect 663 225 664 226
rect 665 225 666 226
rect 460 600 461 601
rect 462 600 463 601
rect 463 600 464 601
rect 465 600 466 601
rect 460 601 466 605
rect 460 605 461 606
rect 462 605 463 606
rect 463 605 464 606
rect 465 605 466 606
rect 580 140 581 141
rect 582 140 583 141
rect 583 140 584 141
rect 585 140 586 141
rect 580 141 586 145
rect 580 145 581 146
rect 582 145 583 146
rect 583 145 584 146
rect 585 145 586 146
rect 60 420 61 421
rect 62 420 63 421
rect 63 420 64 421
rect 65 420 66 421
rect 60 421 66 425
rect 60 425 61 426
rect 62 425 63 426
rect 63 425 64 426
rect 65 425 66 426
rect 460 100 461 101
rect 462 100 463 101
rect 463 100 464 101
rect 465 100 466 101
rect 460 101 466 105
rect 460 105 461 106
rect 462 105 463 106
rect 463 105 464 106
rect 465 105 466 106
rect 560 120 561 121
rect 562 120 563 121
rect 563 120 564 121
rect 565 120 566 121
rect 560 121 566 125
rect 560 125 561 126
rect 562 125 563 126
rect 563 125 564 126
rect 565 125 566 126
rect 540 200 541 201
rect 542 200 543 201
rect 543 200 544 201
rect 545 200 546 201
rect 540 201 546 205
rect 540 205 541 206
rect 542 205 543 206
rect 543 205 544 206
rect 545 205 546 206
rect 420 500 421 501
rect 422 500 423 501
rect 423 500 424 501
rect 425 500 426 501
rect 420 501 426 505
rect 420 505 421 506
rect 422 505 423 506
rect 423 505 424 506
rect 425 505 426 506
rect 300 220 301 221
rect 302 220 303 221
rect 303 220 304 221
rect 305 220 306 221
rect 300 221 306 225
rect 300 225 301 226
rect 302 225 303 226
rect 303 225 304 226
rect 305 225 306 226
rect 540 340 541 341
rect 542 340 543 341
rect 543 340 544 341
rect 545 340 546 341
rect 540 341 546 345
rect 540 345 541 346
rect 542 345 543 346
rect 543 345 544 346
rect 545 345 546 346
rect 240 440 241 441
rect 242 440 243 441
rect 243 440 244 441
rect 245 440 246 441
rect 240 441 246 445
rect 240 445 241 446
rect 242 445 243 446
rect 243 445 244 446
rect 245 445 246 446
rect 480 460 481 461
rect 482 460 483 461
rect 483 460 484 461
rect 485 460 486 461
rect 480 461 486 465
rect 480 465 481 466
rect 482 465 483 466
rect 483 465 484 466
rect 485 465 486 466
rect 260 40 261 41
rect 262 40 263 41
rect 263 40 264 41
rect 265 40 266 41
rect 260 41 266 45
rect 260 45 261 46
rect 262 45 263 46
rect 263 45 264 46
rect 265 45 266 46
rect 560 420 561 421
rect 562 420 563 421
rect 563 420 564 421
rect 565 420 566 421
rect 560 421 566 425
rect 560 425 561 426
rect 562 425 563 426
rect 563 425 564 426
rect 565 425 566 426
rect 340 140 341 141
rect 342 140 343 141
rect 343 140 344 141
rect 345 140 346 141
rect 340 141 346 145
rect 340 145 341 146
rect 342 145 343 146
rect 343 145 344 146
rect 345 145 346 146
rect 600 500 601 501
rect 602 500 603 501
rect 603 500 604 501
rect 605 500 606 501
rect 600 501 606 505
rect 600 505 601 506
rect 602 505 603 506
rect 603 505 604 506
rect 605 505 606 506
rect 100 420 101 421
rect 102 420 103 421
rect 103 420 104 421
rect 105 420 106 421
rect 100 421 106 425
rect 100 425 101 426
rect 102 425 103 426
rect 103 425 104 426
rect 105 425 106 426
rect 520 620 521 621
rect 522 620 523 621
rect 523 620 524 621
rect 525 620 526 621
rect 520 621 526 625
rect 520 625 521 626
rect 522 625 523 626
rect 523 625 524 626
rect 525 625 526 626
rect 640 220 641 221
rect 642 220 643 221
rect 643 220 644 221
rect 645 220 646 221
rect 640 221 646 225
rect 640 225 641 226
rect 642 225 643 226
rect 643 225 644 226
rect 645 225 646 226
rect 300 60 301 61
rect 302 60 303 61
rect 303 60 304 61
rect 305 60 306 61
rect 300 61 306 65
rect 300 65 301 66
rect 302 65 303 66
rect 303 65 304 66
rect 305 65 306 66
rect 240 60 241 61
rect 242 60 243 61
rect 243 60 244 61
rect 245 60 246 61
rect 240 61 246 65
rect 240 65 241 66
rect 242 65 243 66
rect 243 65 244 66
rect 245 65 246 66
rect 360 460 361 461
rect 362 460 363 461
rect 363 460 364 461
rect 365 460 366 461
rect 360 461 366 465
rect 360 465 361 466
rect 362 465 363 466
rect 363 465 364 466
rect 365 465 366 466
rect 400 600 401 601
rect 402 600 403 601
rect 403 600 404 601
rect 405 600 406 601
rect 400 601 406 605
rect 400 605 401 606
rect 402 605 403 606
rect 403 605 404 606
rect 405 605 406 606
rect 500 460 501 461
rect 502 460 503 461
rect 503 460 504 461
rect 505 460 506 461
rect 500 461 506 465
rect 500 465 501 466
rect 502 465 503 466
rect 503 465 504 466
rect 505 465 506 466
rect 240 180 241 181
rect 242 180 243 181
rect 243 180 244 181
rect 245 180 246 181
rect 240 181 246 185
rect 240 185 241 186
rect 242 185 243 186
rect 243 185 244 186
rect 245 185 246 186
rect 420 580 421 581
rect 422 580 423 581
rect 423 580 424 581
rect 425 580 426 581
rect 420 581 426 585
rect 420 585 421 586
rect 422 585 423 586
rect 423 585 424 586
rect 425 585 426 586
rect 200 580 201 581
rect 202 580 203 581
rect 203 580 204 581
rect 205 580 206 581
rect 200 581 206 585
rect 200 585 201 586
rect 202 585 203 586
rect 203 585 204 586
rect 205 585 206 586
rect 300 640 301 641
rect 302 640 303 641
rect 303 640 304 641
rect 305 640 306 641
rect 300 641 306 645
rect 300 645 301 646
rect 302 645 303 646
rect 303 645 304 646
rect 305 645 306 646
rect 240 360 241 361
rect 242 360 243 361
rect 243 360 244 361
rect 245 360 246 361
rect 240 361 246 365
rect 240 365 241 366
rect 242 365 243 366
rect 243 365 244 366
rect 245 365 246 366
rect 500 60 501 61
rect 502 60 503 61
rect 503 60 504 61
rect 505 60 506 61
rect 500 61 506 65
rect 500 65 501 66
rect 502 65 503 66
rect 503 65 504 66
rect 505 65 506 66
rect 460 560 461 561
rect 462 560 463 561
rect 463 560 464 561
rect 465 560 466 561
rect 460 561 466 565
rect 460 565 461 566
rect 462 565 463 566
rect 463 565 464 566
rect 465 565 466 566
rect 420 240 421 241
rect 422 240 423 241
rect 423 240 424 241
rect 425 240 426 241
rect 420 241 426 245
rect 420 245 421 246
rect 422 245 423 246
rect 423 245 424 246
rect 425 245 426 246
rect 340 160 341 161
rect 342 160 343 161
rect 343 160 344 161
rect 345 160 346 161
rect 340 161 346 165
rect 340 165 341 166
rect 342 165 343 166
rect 343 165 344 166
rect 345 165 346 166
rect 580 200 581 201
rect 582 200 583 201
rect 583 200 584 201
rect 585 200 586 201
rect 580 201 586 205
rect 580 205 581 206
rect 582 205 583 206
rect 583 205 584 206
rect 585 205 586 206
rect 140 220 141 221
rect 142 220 143 221
rect 143 220 144 221
rect 145 220 146 221
rect 140 221 146 225
rect 140 225 141 226
rect 142 225 143 226
rect 143 225 144 226
rect 145 225 146 226
rect 340 520 341 521
rect 342 520 343 521
rect 343 520 344 521
rect 345 520 346 521
rect 340 521 346 525
rect 340 525 341 526
rect 342 525 343 526
rect 343 525 344 526
rect 345 525 346 526
rect 120 380 121 381
rect 122 380 123 381
rect 123 380 124 381
rect 125 380 126 381
rect 120 381 126 385
rect 120 385 121 386
rect 122 385 123 386
rect 123 385 124 386
rect 125 385 126 386
rect 620 320 621 321
rect 622 320 623 321
rect 623 320 624 321
rect 625 320 626 321
rect 620 321 626 325
rect 620 325 621 326
rect 622 325 623 326
rect 623 325 624 326
rect 625 325 626 326
rect 120 400 121 401
rect 122 400 123 401
rect 123 400 124 401
rect 125 400 126 401
rect 120 401 126 405
rect 120 405 121 406
rect 122 405 123 406
rect 123 405 124 406
rect 125 405 126 406
rect 660 300 661 301
rect 662 300 663 301
rect 663 300 664 301
rect 665 300 666 301
rect 660 301 666 305
rect 660 305 661 306
rect 662 305 663 306
rect 663 305 664 306
rect 665 305 666 306
rect 480 200 481 201
rect 482 200 483 201
rect 483 200 484 201
rect 485 200 486 201
rect 480 201 486 205
rect 480 205 481 206
rect 482 205 483 206
rect 483 205 484 206
rect 485 205 486 206
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect 140 160 141 161
rect 142 160 143 161
rect 143 160 144 161
rect 145 160 146 161
rect 140 161 146 165
rect 140 165 141 166
rect 142 165 143 166
rect 143 165 144 166
rect 145 165 146 166
rect 60 240 61 241
rect 62 240 63 241
rect 63 240 64 241
rect 65 240 66 241
rect 60 241 66 245
rect 60 245 61 246
rect 62 245 63 246
rect 63 245 64 246
rect 65 245 66 246
rect 420 460 421 461
rect 422 460 423 461
rect 423 460 424 461
rect 425 460 426 461
rect 420 461 426 465
rect 420 465 421 466
rect 422 465 423 466
rect 423 465 424 466
rect 425 465 426 466
rect 220 240 221 241
rect 222 240 223 241
rect 223 240 224 241
rect 225 240 226 241
rect 220 241 226 245
rect 220 245 221 246
rect 222 245 223 246
rect 223 245 224 246
rect 225 245 226 246
rect 260 620 261 621
rect 262 620 263 621
rect 263 620 264 621
rect 265 620 266 621
rect 260 621 266 625
rect 260 625 261 626
rect 262 625 263 626
rect 263 625 264 626
rect 265 625 266 626
rect 240 240 241 241
rect 242 240 243 241
rect 243 240 244 241
rect 245 240 246 241
rect 240 241 246 245
rect 240 245 241 246
rect 242 245 243 246
rect 243 245 244 246
rect 245 245 246 246
rect 80 300 81 301
rect 82 300 83 301
rect 83 300 84 301
rect 85 300 86 301
rect 80 301 86 305
rect 80 305 81 306
rect 82 305 83 306
rect 83 305 84 306
rect 85 305 86 306
rect 160 300 161 301
rect 162 300 163 301
rect 163 300 164 301
rect 165 300 166 301
rect 160 301 166 305
rect 160 305 161 306
rect 162 305 163 306
rect 163 305 164 306
rect 165 305 166 306
rect 40 520 41 521
rect 42 520 43 521
rect 43 520 44 521
rect 45 520 46 521
rect 40 521 46 525
rect 40 525 41 526
rect 42 525 43 526
rect 43 525 44 526
rect 45 525 46 526
rect 520 280 521 281
rect 522 280 523 281
rect 523 280 524 281
rect 525 280 526 281
rect 520 281 526 285
rect 520 285 521 286
rect 522 285 523 286
rect 523 285 524 286
rect 525 285 526 286
rect 580 500 581 501
rect 582 500 583 501
rect 583 500 584 501
rect 585 500 586 501
rect 580 501 586 505
rect 580 505 581 506
rect 582 505 583 506
rect 583 505 584 506
rect 585 505 586 506
rect 100 380 101 381
rect 102 380 103 381
rect 103 380 104 381
rect 105 380 106 381
rect 100 381 106 385
rect 100 385 101 386
rect 102 385 103 386
rect 103 385 104 386
rect 105 385 106 386
rect 220 260 221 261
rect 222 260 223 261
rect 223 260 224 261
rect 225 260 226 261
rect 220 261 226 265
rect 220 265 221 266
rect 222 265 223 266
rect 223 265 224 266
rect 225 265 226 266
rect 100 360 101 361
rect 102 360 103 361
rect 103 360 104 361
rect 105 360 106 361
rect 100 361 106 365
rect 100 365 101 366
rect 102 365 103 366
rect 103 365 104 366
rect 105 365 106 366
rect 80 140 81 141
rect 82 140 83 141
rect 83 140 84 141
rect 85 140 86 141
rect 80 141 86 145
rect 80 145 81 146
rect 82 145 83 146
rect 83 145 84 146
rect 85 145 86 146
rect 40 140 41 141
rect 42 140 43 141
rect 43 140 44 141
rect 45 140 46 141
rect 40 141 46 145
rect 40 145 41 146
rect 42 145 43 146
rect 43 145 44 146
rect 45 145 46 146
rect 340 380 341 381
rect 342 380 343 381
rect 343 380 344 381
rect 345 380 346 381
rect 340 381 346 385
rect 340 385 341 386
rect 342 385 343 386
rect 343 385 344 386
rect 345 385 346 386
rect 280 500 281 501
rect 282 500 283 501
rect 283 500 284 501
rect 285 500 286 501
rect 280 501 286 505
rect 280 505 281 506
rect 282 505 283 506
rect 283 505 284 506
rect 285 505 286 506
rect 640 320 641 321
rect 642 320 643 321
rect 643 320 644 321
rect 645 320 646 321
rect 640 321 646 325
rect 640 325 641 326
rect 642 325 643 326
rect 643 325 644 326
rect 645 325 646 326
rect 440 140 441 141
rect 442 140 443 141
rect 443 140 444 141
rect 445 140 446 141
rect 440 141 446 145
rect 440 145 441 146
rect 442 145 443 146
rect 443 145 444 146
rect 445 145 446 146
rect 280 160 281 161
rect 282 160 283 161
rect 283 160 284 161
rect 285 160 286 161
rect 280 161 286 165
rect 280 165 281 166
rect 282 165 283 166
rect 283 165 284 166
rect 285 165 286 166
rect 140 180 141 181
rect 142 180 143 181
rect 143 180 144 181
rect 145 180 146 181
rect 140 181 146 185
rect 140 185 141 186
rect 142 185 143 186
rect 143 185 144 186
rect 145 185 146 186
rect 360 400 361 401
rect 362 400 363 401
rect 363 400 364 401
rect 365 400 366 401
rect 360 401 366 405
rect 360 405 361 406
rect 362 405 363 406
rect 363 405 364 406
rect 365 405 366 406
rect 0 180 1 181
rect 2 180 3 181
rect 3 180 4 181
rect 5 180 6 181
rect 0 181 6 185
rect 0 185 1 186
rect 2 185 3 186
rect 3 185 4 186
rect 5 185 6 186
rect 480 580 481 581
rect 482 580 483 581
rect 483 580 484 581
rect 485 580 486 581
rect 480 581 486 585
rect 480 585 481 586
rect 482 585 483 586
rect 483 585 484 586
rect 485 585 486 586
rect 200 620 201 621
rect 202 620 203 621
rect 203 620 204 621
rect 205 620 206 621
rect 200 621 206 625
rect 200 625 201 626
rect 202 625 203 626
rect 203 625 204 626
rect 205 625 206 626
rect 160 580 161 581
rect 162 580 163 581
rect 163 580 164 581
rect 165 580 166 581
rect 160 581 166 585
rect 160 585 161 586
rect 162 585 163 586
rect 163 585 164 586
rect 165 585 166 586
rect 180 320 181 321
rect 182 320 183 321
rect 183 320 184 321
rect 185 320 186 321
rect 180 321 186 325
rect 180 325 181 326
rect 182 325 183 326
rect 183 325 184 326
rect 185 325 186 326
rect 60 100 61 101
rect 62 100 63 101
rect 63 100 64 101
rect 65 100 66 101
rect 60 101 66 105
rect 60 105 61 106
rect 62 105 63 106
rect 63 105 64 106
rect 65 105 66 106
rect 220 120 221 121
rect 222 120 223 121
rect 223 120 224 121
rect 225 120 226 121
rect 220 121 226 125
rect 220 125 221 126
rect 222 125 223 126
rect 223 125 224 126
rect 225 125 226 126
<< polysilicon >>
rect 421 439 422 441
rect 424 439 425 441
rect 421 445 422 447
rect 424 445 425 447
rect 361 279 362 281
rect 364 279 365 281
rect 361 285 362 287
rect 364 285 365 287
rect 81 479 82 481
rect 84 479 85 481
rect 81 485 82 487
rect 84 485 85 487
rect 121 159 122 161
rect 124 159 125 161
rect 121 165 122 167
rect 124 165 125 167
rect 461 579 462 581
rect 464 579 465 581
rect 461 585 462 587
rect 464 585 465 587
rect 421 159 422 161
rect 424 159 425 161
rect 421 165 422 167
rect 424 165 425 167
rect 521 19 522 21
rect 524 19 525 21
rect 521 25 522 27
rect 524 25 525 27
rect 481 439 482 441
rect 484 439 485 441
rect 481 445 482 447
rect 484 445 485 447
rect 501 179 502 181
rect 504 179 505 181
rect 501 185 502 187
rect 504 185 505 187
rect 381 99 382 101
rect 384 99 385 101
rect 381 105 382 107
rect 384 105 385 107
rect 581 279 582 281
rect 584 279 585 281
rect 581 285 582 287
rect 584 285 585 287
rect 601 239 602 241
rect 604 239 605 241
rect 601 245 602 247
rect 604 245 605 247
rect 321 159 322 161
rect 324 159 325 161
rect 321 165 322 167
rect 324 165 325 167
rect 341 459 342 461
rect 344 459 345 461
rect 341 465 342 467
rect 344 465 345 467
rect 41 279 42 281
rect 44 279 45 281
rect 41 285 42 287
rect 44 285 45 287
rect 261 499 262 501
rect 264 499 265 501
rect 261 505 262 507
rect 264 505 265 507
rect 481 359 482 361
rect 484 359 485 361
rect 481 365 482 367
rect 484 365 485 367
rect 441 319 442 321
rect 444 319 445 321
rect 441 325 442 327
rect 444 325 445 327
rect 281 59 282 61
rect 284 59 285 61
rect 281 65 282 67
rect 284 65 285 67
rect 541 499 542 501
rect 544 499 545 501
rect 541 505 542 507
rect 544 505 545 507
rect 401 359 402 361
rect 404 359 405 361
rect 401 365 402 367
rect 404 365 405 367
rect 461 139 462 141
rect 464 139 465 141
rect 461 145 462 147
rect 464 145 465 147
rect 301 179 302 181
rect 304 179 305 181
rect 301 185 302 187
rect 304 185 305 187
rect 341 239 342 241
rect 344 239 345 241
rect 341 245 342 247
rect 344 245 345 247
rect 201 39 202 41
rect 204 39 205 41
rect 201 45 202 47
rect 204 45 205 47
rect 261 379 262 381
rect 264 379 265 381
rect 261 385 262 387
rect 264 385 265 387
rect 501 559 502 561
rect 504 559 505 561
rect 501 565 502 567
rect 504 565 505 567
rect 221 159 222 161
rect 224 159 225 161
rect 221 165 222 167
rect 224 165 225 167
rect 281 519 282 521
rect 284 519 285 521
rect 281 525 282 527
rect 284 525 285 527
rect 201 479 202 481
rect 204 479 205 481
rect 201 485 202 487
rect 204 485 205 487
rect 461 59 462 61
rect 464 59 465 61
rect 461 65 462 67
rect 464 65 465 67
rect 181 459 182 461
rect 184 459 185 461
rect 181 465 182 467
rect 184 465 185 467
rect 321 19 322 21
rect 324 19 325 21
rect 321 25 322 27
rect 324 25 325 27
rect 321 279 322 281
rect 324 279 325 281
rect 321 285 322 287
rect 324 285 325 287
rect 561 259 562 261
rect 564 259 565 261
rect 561 265 562 267
rect 564 265 565 267
rect 561 319 562 321
rect 564 319 565 321
rect 561 325 562 327
rect 564 325 565 327
rect 661 359 662 361
rect 664 359 665 361
rect 661 365 662 367
rect 664 365 665 367
rect 341 99 342 101
rect 344 99 345 101
rect 341 105 342 107
rect 344 105 345 107
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect 381 139 382 141
rect 384 139 385 141
rect 381 145 382 147
rect 384 145 385 147
rect 141 379 142 381
rect 144 379 145 381
rect 141 385 142 387
rect 144 385 145 387
rect 321 -1 322 1
rect 324 -1 325 1
rect 321 5 322 7
rect 324 5 325 7
rect 341 399 342 401
rect 344 399 345 401
rect 341 405 342 407
rect 344 405 345 407
rect 481 399 482 401
rect 484 399 485 401
rect 481 405 482 407
rect 484 405 485 407
rect 161 519 162 521
rect 164 519 165 521
rect 161 525 162 527
rect 164 525 165 527
rect 281 379 282 381
rect 284 379 285 381
rect 281 385 282 387
rect 284 385 285 387
rect 421 419 422 421
rect 424 419 425 421
rect 421 425 422 427
rect 424 425 425 427
rect 541 539 542 541
rect 544 539 545 541
rect 541 545 542 547
rect 544 545 545 547
rect 141 519 142 521
rect 144 519 145 521
rect 141 525 142 527
rect 144 525 145 527
rect 461 199 462 201
rect 464 199 465 201
rect 461 205 462 207
rect 464 205 465 207
rect 381 539 382 541
rect 384 539 385 541
rect 381 545 382 547
rect 384 545 385 547
rect 461 179 462 181
rect 464 179 465 181
rect 461 185 462 187
rect 464 185 465 187
rect 61 399 62 401
rect 64 399 65 401
rect 61 405 62 407
rect 64 405 65 407
rect 241 139 242 141
rect 244 139 245 141
rect 241 145 242 147
rect 244 145 245 147
rect 21 279 22 281
rect 24 279 25 281
rect 21 285 22 287
rect 24 285 25 287
rect 481 599 482 601
rect 484 599 485 601
rect 481 605 482 607
rect 484 605 485 607
rect 381 359 382 361
rect 384 359 385 361
rect 381 365 382 367
rect 384 365 385 367
rect 241 119 242 121
rect 244 119 245 121
rect 241 125 242 127
rect 244 125 245 127
rect 421 639 422 641
rect 424 639 425 641
rect 421 645 422 647
rect 424 645 425 647
rect 601 159 602 161
rect 604 159 605 161
rect 601 165 602 167
rect 604 165 605 167
rect 381 659 382 661
rect 384 659 385 661
rect 381 665 382 667
rect 384 665 385 667
rect 281 119 282 121
rect 284 119 285 121
rect 281 125 282 127
rect 284 125 285 127
rect 301 439 302 441
rect 304 439 305 441
rect 301 445 302 447
rect 304 445 305 447
rect 281 539 282 541
rect 284 539 285 541
rect 281 545 282 547
rect 284 545 285 547
rect 201 79 202 81
rect 204 79 205 81
rect 201 85 202 87
rect 204 85 205 87
rect 21 179 22 181
rect 24 179 25 181
rect 21 185 22 187
rect 24 185 25 187
rect 401 99 402 101
rect 404 99 405 101
rect 401 105 402 107
rect 404 105 405 107
rect 481 639 482 641
rect 484 639 485 641
rect 481 645 482 647
rect 484 645 485 647
rect 361 519 362 521
rect 364 519 365 521
rect 361 525 362 527
rect 364 525 365 527
rect 81 119 82 121
rect 84 119 85 121
rect 81 125 82 127
rect 84 125 85 127
rect 321 119 322 121
rect 324 119 325 121
rect 321 125 322 127
rect 324 125 325 127
rect 301 199 302 201
rect 304 199 305 201
rect 301 205 302 207
rect 304 205 305 207
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect 301 479 302 481
rect 304 479 305 481
rect 301 485 302 487
rect 304 485 305 487
rect 41 339 42 341
rect 44 339 45 341
rect 41 345 42 347
rect 44 345 45 347
rect 481 239 482 241
rect 484 239 485 241
rect 481 245 482 247
rect 484 245 485 247
rect 201 259 202 261
rect 204 259 205 261
rect 201 265 202 267
rect 204 265 205 267
rect 381 439 382 441
rect 384 439 385 441
rect 381 445 382 447
rect 384 445 385 447
rect 281 299 282 301
rect 284 299 285 301
rect 281 305 282 307
rect 284 305 285 307
rect 621 199 622 201
rect 624 199 625 201
rect 621 205 622 207
rect 624 205 625 207
rect 321 479 322 481
rect 324 479 325 481
rect 321 485 322 487
rect 324 485 325 487
rect 601 519 602 521
rect 604 519 605 521
rect 601 525 602 527
rect 604 525 605 527
rect 121 619 122 621
rect 124 619 125 621
rect 121 625 122 627
rect 124 625 125 627
rect 401 199 402 201
rect 404 199 405 201
rect 401 205 402 207
rect 404 205 405 207
rect 21 399 22 401
rect 24 399 25 401
rect 21 405 22 407
rect 24 405 25 407
rect 281 -1 282 1
rect 284 -1 285 1
rect 281 5 282 7
rect 284 5 285 7
rect 281 399 282 401
rect 284 399 285 401
rect 281 405 282 407
rect 284 405 285 407
rect 461 239 462 241
rect 464 239 465 241
rect 461 245 462 247
rect 464 245 465 247
rect 301 279 302 281
rect 304 279 305 281
rect 301 285 302 287
rect 304 285 305 287
rect 441 599 442 601
rect 444 599 445 601
rect 441 605 442 607
rect 444 605 445 607
rect 121 419 122 421
rect 124 419 125 421
rect 121 425 122 427
rect 124 425 125 427
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect 101 539 102 541
rect 104 539 105 541
rect 101 545 102 547
rect 104 545 105 547
rect 341 79 342 81
rect 344 79 345 81
rect 341 85 342 87
rect 344 85 345 87
rect 221 439 222 441
rect 224 439 225 441
rect 221 445 222 447
rect 224 445 225 447
rect 341 179 342 181
rect 344 179 345 181
rect 341 185 342 187
rect 344 185 345 187
rect 361 319 362 321
rect 364 319 365 321
rect 361 325 362 327
rect 364 325 365 327
rect 41 239 42 241
rect 44 239 45 241
rect 41 245 42 247
rect 44 245 45 247
rect 181 659 182 661
rect 184 659 185 661
rect 181 665 182 667
rect 184 665 185 667
rect 521 39 522 41
rect 524 39 525 41
rect 521 45 522 47
rect 524 45 525 47
rect 241 299 242 301
rect 244 299 245 301
rect 241 305 242 307
rect 244 305 245 307
rect 361 159 362 161
rect 364 159 365 161
rect 361 165 362 167
rect 364 165 365 167
rect 401 519 402 521
rect 404 519 405 521
rect 401 525 402 527
rect 404 525 405 527
rect 341 639 342 641
rect 344 639 345 641
rect 341 645 342 647
rect 344 645 345 647
rect 201 159 202 161
rect 204 159 205 161
rect 201 165 202 167
rect 204 165 205 167
rect 21 99 22 101
rect 24 99 25 101
rect 21 105 22 107
rect 24 105 25 107
rect 341 479 342 481
rect 344 479 345 481
rect 341 485 342 487
rect 344 485 345 487
rect 161 259 162 261
rect 164 259 165 261
rect 161 265 162 267
rect 164 265 165 267
rect 501 139 502 141
rect 504 139 505 141
rect 501 145 502 147
rect 504 145 505 147
rect 401 39 402 41
rect 404 39 405 41
rect 401 45 402 47
rect 404 45 405 47
rect 241 539 242 541
rect 244 539 245 541
rect 241 545 242 547
rect 244 545 245 547
rect 521 539 522 541
rect 524 539 525 541
rect 521 545 522 547
rect 524 545 525 547
rect 341 319 342 321
rect 344 319 345 321
rect 341 325 342 327
rect 344 325 345 327
rect 381 459 382 461
rect 384 459 385 461
rect 381 465 382 467
rect 384 465 385 467
rect 101 219 102 221
rect 104 219 105 221
rect 101 225 102 227
rect 104 225 105 227
rect 601 179 602 181
rect 604 179 605 181
rect 601 185 602 187
rect 604 185 605 187
rect 461 339 462 341
rect 464 339 465 341
rect 461 345 462 347
rect 464 345 465 347
rect 81 159 82 161
rect 84 159 85 161
rect 81 165 82 167
rect 84 165 85 167
rect 521 199 522 201
rect 524 199 525 201
rect 521 205 522 207
rect 524 205 525 207
rect 201 359 202 361
rect 204 359 205 361
rect 201 365 202 367
rect 204 365 205 367
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect 121 139 122 141
rect 124 139 125 141
rect 121 145 122 147
rect 124 145 125 147
rect 161 419 162 421
rect 164 419 165 421
rect 161 425 162 427
rect 164 425 165 427
rect 321 399 322 401
rect 324 399 325 401
rect 321 405 322 407
rect 324 405 325 407
rect 461 519 462 521
rect 464 519 465 521
rect 461 525 462 527
rect 464 525 465 527
rect 361 379 362 381
rect 364 379 365 381
rect 361 385 362 387
rect 364 385 365 387
rect 261 439 262 441
rect 264 439 265 441
rect 261 445 262 447
rect 264 445 265 447
rect 281 439 282 441
rect 284 439 285 441
rect 281 445 282 447
rect 284 445 285 447
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect 501 379 502 381
rect 504 379 505 381
rect 501 385 502 387
rect 504 385 505 387
rect 501 339 502 341
rect 504 339 505 341
rect 501 345 502 347
rect 504 345 505 347
rect 341 539 342 541
rect 344 539 345 541
rect 341 545 342 547
rect 344 545 345 547
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect 541 379 542 381
rect 544 379 545 381
rect 541 385 542 387
rect 544 385 545 387
rect 261 259 262 261
rect 264 259 265 261
rect 261 265 262 267
rect 264 265 265 267
rect 441 219 442 221
rect 444 219 445 221
rect 441 225 442 227
rect 444 225 445 227
rect 161 239 162 241
rect 164 239 165 241
rect 161 245 162 247
rect 164 245 165 247
rect 481 539 482 541
rect 484 539 485 541
rect 481 545 482 547
rect 484 545 485 547
rect 381 559 382 561
rect 384 559 385 561
rect 381 565 382 567
rect 384 565 385 567
rect 441 399 442 401
rect 444 399 445 401
rect 441 405 442 407
rect 444 405 445 407
rect 621 179 622 181
rect 624 179 625 181
rect 621 185 622 187
rect 624 185 625 187
rect 301 299 302 301
rect 304 299 305 301
rect 301 305 302 307
rect 304 305 305 307
rect 541 599 542 601
rect 544 599 545 601
rect 541 605 542 607
rect 544 605 545 607
rect 21 239 22 241
rect 24 239 25 241
rect 21 245 22 247
rect 24 245 25 247
rect 321 539 322 541
rect 324 539 325 541
rect 321 545 322 547
rect 324 545 325 547
rect 361 659 362 661
rect 364 659 365 661
rect 361 665 362 667
rect 364 665 365 667
rect 281 339 282 341
rect 284 339 285 341
rect 281 345 282 347
rect 284 345 285 347
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect 441 459 442 461
rect 444 459 445 461
rect 441 465 442 467
rect 444 465 445 467
rect 261 139 262 141
rect 264 139 265 141
rect 261 145 262 147
rect 264 145 265 147
rect 581 239 582 241
rect 584 239 585 241
rect 581 245 582 247
rect 584 245 585 247
rect 221 59 222 61
rect 224 59 225 61
rect 221 65 222 67
rect 224 65 225 67
rect 401 539 402 541
rect 404 539 405 541
rect 401 545 402 547
rect 404 545 405 547
rect 281 419 282 421
rect 284 419 285 421
rect 281 425 282 427
rect 284 425 285 427
rect 321 499 322 501
rect 324 499 325 501
rect 321 505 322 507
rect 324 505 325 507
rect 321 459 322 461
rect 324 459 325 461
rect 321 465 322 467
rect 324 465 325 467
rect 1 259 2 261
rect 4 259 5 261
rect 1 265 2 267
rect 4 265 5 267
rect 241 459 242 461
rect 244 459 245 461
rect 241 465 242 467
rect 244 465 245 467
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect 141 119 142 121
rect 144 119 145 121
rect 141 125 142 127
rect 144 125 145 127
rect 561 179 562 181
rect 564 179 565 181
rect 561 185 562 187
rect 564 185 565 187
rect 61 159 62 161
rect 64 159 65 161
rect 61 165 62 167
rect 64 165 65 167
rect 521 139 522 141
rect 524 139 525 141
rect 521 145 522 147
rect 524 145 525 147
rect 261 339 262 341
rect 264 339 265 341
rect 261 345 262 347
rect 264 345 265 347
rect 321 219 322 221
rect 324 219 325 221
rect 321 225 322 227
rect 324 225 325 227
rect 441 439 442 441
rect 444 439 445 441
rect 441 445 442 447
rect 444 445 445 447
rect 201 639 202 641
rect 204 639 205 641
rect 201 645 202 647
rect 204 645 205 647
rect 361 499 362 501
rect 364 499 365 501
rect 361 505 362 507
rect 364 505 365 507
rect 21 499 22 501
rect 24 499 25 501
rect 21 505 22 507
rect 24 505 25 507
rect 381 59 382 61
rect 384 59 385 61
rect 381 65 382 67
rect 384 65 385 67
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect 341 219 342 221
rect 344 219 345 221
rect 341 225 342 227
rect 344 225 345 227
rect 461 379 462 381
rect 464 379 465 381
rect 461 385 462 387
rect 464 385 465 387
rect 661 279 662 281
rect 664 279 665 281
rect 661 285 662 287
rect 664 285 665 287
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect 41 259 42 261
rect 44 259 45 261
rect 41 265 42 267
rect 44 265 45 267
rect 241 479 242 481
rect 244 479 245 481
rect 241 485 242 487
rect 244 485 245 487
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect 661 339 662 341
rect 664 339 665 341
rect 661 345 662 347
rect 664 345 665 347
rect 141 439 142 441
rect 144 439 145 441
rect 141 445 142 447
rect 144 445 145 447
rect 521 99 522 101
rect 524 99 525 101
rect 521 105 522 107
rect 524 105 525 107
rect 621 399 622 401
rect 624 399 625 401
rect 621 405 622 407
rect 624 405 625 407
rect 281 319 282 321
rect 284 319 285 321
rect 281 325 282 327
rect 284 325 285 327
rect 61 119 62 121
rect 64 119 65 121
rect 61 125 62 127
rect 64 125 65 127
rect 341 119 342 121
rect 344 119 345 121
rect 341 125 342 127
rect 344 125 345 127
rect 441 339 442 341
rect 444 339 445 341
rect 441 345 442 347
rect 444 345 445 347
rect 521 359 522 361
rect 524 359 525 361
rect 521 365 522 367
rect 524 365 525 367
rect 321 379 322 381
rect 324 379 325 381
rect 321 385 322 387
rect 324 385 325 387
rect 601 399 602 401
rect 604 399 605 401
rect 601 405 602 407
rect 604 405 605 407
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect 601 259 602 261
rect 604 259 605 261
rect 601 265 602 267
rect 604 265 605 267
rect 221 39 222 41
rect 224 39 225 41
rect 221 45 222 47
rect 224 45 225 47
rect 121 119 122 121
rect 124 119 125 121
rect 121 125 122 127
rect 124 125 125 127
rect 501 499 502 501
rect 504 499 505 501
rect 501 505 502 507
rect 504 505 505 507
rect 141 499 142 501
rect 144 499 145 501
rect 141 505 142 507
rect 144 505 145 507
rect 441 659 442 661
rect 444 659 445 661
rect 441 665 442 667
rect 444 665 445 667
rect 401 339 402 341
rect 404 339 405 341
rect 401 345 402 347
rect 404 345 405 347
rect 401 219 402 221
rect 404 219 405 221
rect 401 225 402 227
rect 404 225 405 227
rect 121 319 122 321
rect 124 319 125 321
rect 121 325 122 327
rect 124 325 125 327
rect 421 279 422 281
rect 424 279 425 281
rect 421 285 422 287
rect 424 285 425 287
rect 541 219 542 221
rect 544 219 545 221
rect 541 225 542 227
rect 544 225 545 227
rect 221 179 222 181
rect 224 179 225 181
rect 221 185 222 187
rect 224 185 225 187
rect 281 19 282 21
rect 284 19 285 21
rect 281 25 282 27
rect 284 25 285 27
rect 421 599 422 601
rect 424 599 425 601
rect 421 605 422 607
rect 424 605 425 607
rect 181 119 182 121
rect 184 119 185 121
rect 181 125 182 127
rect 184 125 185 127
rect 461 499 462 501
rect 464 499 465 501
rect 461 505 462 507
rect 464 505 465 507
rect 241 379 242 381
rect 244 379 245 381
rect 241 385 242 387
rect 244 385 245 387
rect 241 219 242 221
rect 244 219 245 221
rect 241 225 242 227
rect 244 225 245 227
rect 301 339 302 341
rect 304 339 305 341
rect 301 345 302 347
rect 304 345 305 347
rect 461 259 462 261
rect 464 259 465 261
rect 461 265 462 267
rect 464 265 465 267
rect 121 439 122 441
rect 124 439 125 441
rect 121 445 122 447
rect 124 445 125 447
rect 181 539 182 541
rect 184 539 185 541
rect 181 545 182 547
rect 184 545 185 547
rect 461 79 462 81
rect 464 79 465 81
rect 461 85 462 87
rect 464 85 465 87
rect 581 299 582 301
rect 584 299 585 301
rect 581 305 582 307
rect 584 305 585 307
rect 461 419 462 421
rect 464 419 465 421
rect 461 425 462 427
rect 464 425 465 427
rect 121 339 122 341
rect 124 339 125 341
rect 121 345 122 347
rect 124 345 125 347
rect 221 319 222 321
rect 224 319 225 321
rect 221 325 222 327
rect 224 325 225 327
rect 421 79 422 81
rect 424 79 425 81
rect 421 85 422 87
rect 424 85 425 87
rect 61 559 62 561
rect 64 559 65 561
rect 61 565 62 567
rect 64 565 65 567
rect 421 219 422 221
rect 424 219 425 221
rect 421 225 422 227
rect 424 225 425 227
rect 321 519 322 521
rect 324 519 325 521
rect 321 525 322 527
rect 324 525 325 527
rect 401 139 402 141
rect 404 139 405 141
rect 401 145 402 147
rect 404 145 405 147
rect 401 119 402 121
rect 404 119 405 121
rect 401 125 402 127
rect 404 125 405 127
rect 381 479 382 481
rect 384 479 385 481
rect 381 485 382 487
rect 384 485 385 487
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect 121 99 122 101
rect 124 99 125 101
rect 121 105 122 107
rect 124 105 125 107
rect 501 99 502 101
rect 504 99 505 101
rect 501 105 502 107
rect 504 105 505 107
rect 301 379 302 381
rect 304 379 305 381
rect 301 385 302 387
rect 304 385 305 387
rect 81 439 82 441
rect 84 439 85 441
rect 81 445 82 447
rect 84 445 85 447
rect 381 599 382 601
rect 384 599 385 601
rect 381 605 382 607
rect 384 605 385 607
rect 201 -1 202 1
rect 204 -1 205 1
rect 201 5 202 7
rect 204 5 205 7
rect 481 339 482 341
rect 484 339 485 341
rect 481 345 482 347
rect 484 345 485 347
rect 221 99 222 101
rect 224 99 225 101
rect 221 105 222 107
rect 224 105 225 107
rect 161 159 162 161
rect 164 159 165 161
rect 161 165 162 167
rect 164 165 165 167
rect 141 259 142 261
rect 144 259 145 261
rect 141 265 142 267
rect 144 265 145 267
rect 101 499 102 501
rect 104 499 105 501
rect 101 505 102 507
rect 104 505 105 507
rect 161 439 162 441
rect 164 439 165 441
rect 161 445 162 447
rect 164 445 165 447
rect 521 579 522 581
rect 524 579 525 581
rect 521 585 522 587
rect 524 585 525 587
rect 301 539 302 541
rect 304 539 305 541
rect 301 545 302 547
rect 304 545 305 547
rect 381 579 382 581
rect 384 579 385 581
rect 381 585 382 587
rect 384 585 385 587
rect 361 179 362 181
rect 364 179 365 181
rect 361 185 362 187
rect 364 185 365 187
rect 21 219 22 221
rect 24 219 25 221
rect 21 225 22 227
rect 24 225 25 227
rect 661 319 662 321
rect 664 319 665 321
rect 661 325 662 327
rect 664 325 665 327
rect 321 79 322 81
rect 324 79 325 81
rect 321 85 322 87
rect 324 85 325 87
rect 321 59 322 61
rect 324 59 325 61
rect 321 65 322 67
rect 324 65 325 67
rect 261 579 262 581
rect 264 579 265 581
rect 261 585 262 587
rect 264 585 265 587
rect 261 59 262 61
rect 264 59 265 61
rect 261 65 262 67
rect 264 65 265 67
rect 221 499 222 501
rect 224 499 225 501
rect 221 505 222 507
rect 224 505 225 507
rect 461 19 462 21
rect 464 19 465 21
rect 461 25 462 27
rect 464 25 465 27
rect 101 399 102 401
rect 104 399 105 401
rect 101 405 102 407
rect 104 405 105 407
rect 381 19 382 21
rect 384 19 385 21
rect 381 25 382 27
rect 384 25 385 27
rect 261 119 262 121
rect 264 119 265 121
rect 261 125 262 127
rect 264 125 265 127
rect 161 179 162 181
rect 164 179 165 181
rect 161 185 162 187
rect 164 185 165 187
rect 341 199 342 201
rect 344 199 345 201
rect 341 205 342 207
rect 344 205 345 207
rect 501 79 502 81
rect 504 79 505 81
rect 501 85 502 87
rect 504 85 505 87
rect 501 359 502 361
rect 504 359 505 361
rect 501 365 502 367
rect 504 365 505 367
rect 581 179 582 181
rect 584 179 585 181
rect 581 185 582 187
rect 584 185 585 187
rect 361 -1 362 1
rect 364 -1 365 1
rect 361 5 362 7
rect 364 5 365 7
rect 521 179 522 181
rect 524 179 525 181
rect 521 185 522 187
rect 524 185 525 187
rect 501 119 502 121
rect 504 119 505 121
rect 501 125 502 127
rect 504 125 505 127
rect 601 299 602 301
rect 604 299 605 301
rect 601 305 602 307
rect 604 305 605 307
rect 101 519 102 521
rect 104 519 105 521
rect 101 525 102 527
rect 104 525 105 527
rect 101 239 102 241
rect 104 239 105 241
rect 101 245 102 247
rect 104 245 105 247
rect 81 179 82 181
rect 84 179 85 181
rect 81 185 82 187
rect 84 185 85 187
rect 261 419 262 421
rect 264 419 265 421
rect 261 425 262 427
rect 264 425 265 427
rect 321 639 322 641
rect 324 639 325 641
rect 321 645 322 647
rect 324 645 325 647
rect 221 599 222 601
rect 224 599 225 601
rect 221 605 222 607
rect 224 605 225 607
rect 501 239 502 241
rect 504 239 505 241
rect 501 245 502 247
rect 504 245 505 247
rect 101 459 102 461
rect 104 459 105 461
rect 101 465 102 467
rect 104 465 105 467
rect 401 379 402 381
rect 404 379 405 381
rect 401 385 402 387
rect 404 385 405 387
rect 201 199 202 201
rect 204 199 205 201
rect 201 205 202 207
rect 204 205 205 207
rect 301 399 302 401
rect 304 399 305 401
rect 301 405 302 407
rect 304 405 305 407
rect 81 559 82 561
rect 84 559 85 561
rect 81 565 82 567
rect 84 565 85 567
rect 241 259 242 261
rect 244 259 245 261
rect 241 265 242 267
rect 244 265 245 267
rect 601 139 602 141
rect 604 139 605 141
rect 601 145 602 147
rect 604 145 605 147
rect 181 19 182 21
rect 184 19 185 21
rect 181 25 182 27
rect 184 25 185 27
rect 601 119 602 121
rect 604 119 605 121
rect 601 125 602 127
rect 604 125 605 127
rect 81 459 82 461
rect 84 459 85 461
rect 81 465 82 467
rect 84 465 85 467
rect 541 279 542 281
rect 544 279 545 281
rect 541 285 542 287
rect 544 285 545 287
rect 201 119 202 121
rect 204 119 205 121
rect 201 125 202 127
rect 204 125 205 127
rect 41 479 42 481
rect 44 479 45 481
rect 41 485 42 487
rect 44 485 45 487
rect 121 539 122 541
rect 124 539 125 541
rect 121 545 122 547
rect 124 545 125 547
rect 421 659 422 661
rect 424 659 425 661
rect 421 665 422 667
rect 424 665 425 667
rect 501 419 502 421
rect 504 419 505 421
rect 501 425 502 427
rect 504 425 505 427
rect 21 299 22 301
rect 24 299 25 301
rect 21 305 22 307
rect 24 305 25 307
rect 581 479 582 481
rect 584 479 585 481
rect 581 485 582 487
rect 584 485 585 487
rect 141 79 142 81
rect 144 79 145 81
rect 141 85 142 87
rect 144 85 145 87
rect 321 179 322 181
rect 324 179 325 181
rect 321 185 322 187
rect 324 185 325 187
rect 21 379 22 381
rect 24 379 25 381
rect 21 385 22 387
rect 24 385 25 387
rect 41 419 42 421
rect 44 419 45 421
rect 41 425 42 427
rect 44 425 45 427
rect 641 359 642 361
rect 644 359 645 361
rect 641 365 642 367
rect 644 365 645 367
rect 401 79 402 81
rect 404 79 405 81
rect 401 85 402 87
rect 404 85 405 87
rect 1 239 2 241
rect 4 239 5 241
rect 1 245 2 247
rect 4 245 5 247
rect 181 239 182 241
rect 184 239 185 241
rect 181 245 182 247
rect 184 245 185 247
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect 281 459 282 461
rect 284 459 285 461
rect 281 465 282 467
rect 284 465 285 467
rect 641 259 642 261
rect 644 259 645 261
rect 641 265 642 267
rect 644 265 645 267
rect 561 219 562 221
rect 564 219 565 221
rect 561 225 562 227
rect 564 225 565 227
rect 441 59 442 61
rect 444 59 445 61
rect 441 65 442 67
rect 444 65 445 67
rect 521 479 522 481
rect 524 479 525 481
rect 521 485 522 487
rect 524 485 525 487
rect 261 99 262 101
rect 264 99 265 101
rect 261 105 262 107
rect 264 105 265 107
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect 261 479 262 481
rect 264 479 265 481
rect 261 485 262 487
rect 264 485 265 487
rect 181 519 182 521
rect 184 519 185 521
rect 181 525 182 527
rect 184 525 185 527
rect 361 259 362 261
rect 364 259 365 261
rect 361 265 362 267
rect 364 265 365 267
rect 321 439 322 441
rect 324 439 325 441
rect 321 445 322 447
rect 324 445 325 447
rect 361 479 362 481
rect 364 479 365 481
rect 361 485 362 487
rect 364 485 365 487
rect 261 159 262 161
rect 264 159 265 161
rect 261 165 262 167
rect 264 165 265 167
rect 661 239 662 241
rect 664 239 665 241
rect 661 245 662 247
rect 664 245 665 247
rect 201 239 202 241
rect 204 239 205 241
rect 201 245 202 247
rect 204 245 205 247
rect 481 319 482 321
rect 484 319 485 321
rect 481 325 482 327
rect 484 325 485 327
rect 121 499 122 501
rect 124 499 125 501
rect 121 505 122 507
rect 124 505 125 507
rect 41 399 42 401
rect 44 399 45 401
rect 41 405 42 407
rect 44 405 45 407
rect 221 279 222 281
rect 224 279 225 281
rect 221 285 222 287
rect 224 285 225 287
rect 281 659 282 661
rect 284 659 285 661
rect 281 665 282 667
rect 284 665 285 667
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect 621 339 622 341
rect 624 339 625 341
rect 621 345 622 347
rect 624 345 625 347
rect 481 619 482 621
rect 484 619 485 621
rect 481 625 482 627
rect 484 625 485 627
rect 181 479 182 481
rect 184 479 185 481
rect 181 485 182 487
rect 184 485 185 487
rect 641 299 642 301
rect 644 299 645 301
rect 641 305 642 307
rect 644 305 645 307
rect 101 479 102 481
rect 104 479 105 481
rect 101 485 102 487
rect 104 485 105 487
rect 501 299 502 301
rect 504 299 505 301
rect 501 305 502 307
rect 504 305 505 307
rect 181 559 182 561
rect 184 559 185 561
rect 181 565 182 567
rect 184 565 185 567
rect 361 299 362 301
rect 364 299 365 301
rect 361 305 362 307
rect 364 305 365 307
rect 261 239 262 241
rect 264 239 265 241
rect 261 245 262 247
rect 264 245 265 247
rect 41 459 42 461
rect 44 459 45 461
rect 41 465 42 467
rect 44 465 45 467
rect 401 579 402 581
rect 404 579 405 581
rect 401 585 402 587
rect 404 585 405 587
rect 201 399 202 401
rect 204 399 205 401
rect 201 405 202 407
rect 204 405 205 407
rect 641 479 642 481
rect 644 479 645 481
rect 641 485 642 487
rect 644 485 645 487
rect 101 99 102 101
rect 104 99 105 101
rect 101 105 102 107
rect 104 105 105 107
rect 401 419 402 421
rect 404 419 405 421
rect 401 425 402 427
rect 404 425 405 427
rect 521 299 522 301
rect 524 299 525 301
rect 521 305 522 307
rect 524 305 525 307
rect 241 319 242 321
rect 244 319 245 321
rect 241 325 242 327
rect 244 325 245 327
rect 281 559 282 561
rect 284 559 285 561
rect 281 565 282 567
rect 284 565 285 567
rect 41 439 42 441
rect 44 439 45 441
rect 41 445 42 447
rect 44 445 45 447
rect 1 159 2 161
rect 4 159 5 161
rect 1 165 2 167
rect 4 165 5 167
rect 261 179 262 181
rect 264 179 265 181
rect 261 185 262 187
rect 264 185 265 187
rect 401 459 402 461
rect 404 459 405 461
rect 401 465 402 467
rect 404 465 405 467
rect 601 379 602 381
rect 604 379 605 381
rect 601 385 602 387
rect 604 385 605 387
rect 161 219 162 221
rect 164 219 165 221
rect 161 225 162 227
rect 164 225 165 227
rect 221 559 222 561
rect 224 559 225 561
rect 221 565 222 567
rect 224 565 225 567
rect 481 159 482 161
rect 484 159 485 161
rect 481 165 482 167
rect 484 165 485 167
rect 301 499 302 501
rect 304 499 305 501
rect 301 505 302 507
rect 304 505 305 507
rect 81 399 82 401
rect 84 399 85 401
rect 81 405 82 407
rect 84 405 85 407
rect 341 339 342 341
rect 344 339 345 341
rect 341 345 342 347
rect 344 345 345 347
rect 401 -1 402 1
rect 404 -1 405 1
rect 401 5 402 7
rect 404 5 405 7
rect 481 179 482 181
rect 484 179 485 181
rect 481 185 482 187
rect 484 185 485 187
rect 421 399 422 401
rect 424 399 425 401
rect 421 405 422 407
rect 424 405 425 407
rect 281 579 282 581
rect 284 579 285 581
rect 281 585 282 587
rect 284 585 285 587
rect 441 119 442 121
rect 444 119 445 121
rect 441 125 442 127
rect 444 125 445 127
rect 181 59 182 61
rect 184 59 185 61
rect 181 65 182 67
rect 184 65 185 67
rect 461 399 462 401
rect 464 399 465 401
rect 461 405 462 407
rect 464 405 465 407
rect 561 399 562 401
rect 564 399 565 401
rect 561 405 562 407
rect 564 405 565 407
rect 541 139 542 141
rect 544 139 545 141
rect 541 145 542 147
rect 544 145 545 147
rect 181 379 182 381
rect 184 379 185 381
rect 181 385 182 387
rect 184 385 185 387
rect 601 439 602 441
rect 604 439 605 441
rect 601 445 602 447
rect 604 445 605 447
rect 481 99 482 101
rect 484 99 485 101
rect 481 105 482 107
rect 484 105 485 107
rect 241 519 242 521
rect 244 519 245 521
rect 241 525 242 527
rect 244 525 245 527
rect 241 579 242 581
rect 244 579 245 581
rect 241 585 242 587
rect 244 585 245 587
rect 381 179 382 181
rect 384 179 385 181
rect 381 185 382 187
rect 384 185 385 187
rect 641 379 642 381
rect 644 379 645 381
rect 641 385 642 387
rect 644 385 645 387
rect 341 499 342 501
rect 344 499 345 501
rect 341 505 342 507
rect 344 505 345 507
rect 61 499 62 501
rect 64 499 65 501
rect 61 505 62 507
rect 64 505 65 507
rect 201 319 202 321
rect 204 319 205 321
rect 201 325 202 327
rect 204 325 205 327
rect 581 159 582 161
rect 584 159 585 161
rect 581 165 582 167
rect 584 165 585 167
rect 121 79 122 81
rect 124 79 125 81
rect 121 85 122 87
rect 124 85 125 87
rect 441 539 442 541
rect 444 539 445 541
rect 441 545 442 547
rect 444 545 445 547
rect 141 59 142 61
rect 144 59 145 61
rect 141 65 142 67
rect 144 65 145 67
rect 1 459 2 461
rect 4 459 5 461
rect 1 465 2 467
rect 4 465 5 467
rect 621 279 622 281
rect 624 279 625 281
rect 621 285 622 287
rect 624 285 625 287
rect 481 559 482 561
rect 484 559 485 561
rect 481 565 482 567
rect 484 565 485 567
rect 21 459 22 461
rect 24 459 25 461
rect 21 465 22 467
rect 24 465 25 467
rect 481 259 482 261
rect 484 259 485 261
rect 481 265 482 267
rect 484 265 485 267
rect 261 539 262 541
rect 264 539 265 541
rect 261 545 262 547
rect 264 545 265 547
rect 261 -1 262 1
rect 264 -1 265 1
rect 261 5 262 7
rect 264 5 265 7
rect 81 259 82 261
rect 84 259 85 261
rect 81 265 82 267
rect 84 265 85 267
rect 481 479 482 481
rect 484 479 485 481
rect 481 485 482 487
rect 484 485 485 487
rect 281 239 282 241
rect 284 239 285 241
rect 281 245 282 247
rect 284 245 285 247
rect 461 639 462 641
rect 464 639 465 641
rect 461 645 462 647
rect 464 645 465 647
rect 461 459 462 461
rect 464 459 465 461
rect 461 465 462 467
rect 464 465 465 467
rect 341 359 342 361
rect 344 359 345 361
rect 341 365 342 367
rect 344 365 345 367
rect 301 139 302 141
rect 304 139 305 141
rect 301 145 302 147
rect 304 145 305 147
rect 661 259 662 261
rect 664 259 665 261
rect 661 265 662 267
rect 664 265 665 267
rect 381 259 382 261
rect 384 259 385 261
rect 381 265 382 267
rect 384 265 385 267
rect 81 59 82 61
rect 84 59 85 61
rect 81 65 82 67
rect 84 65 85 67
rect 341 299 342 301
rect 344 299 345 301
rect 341 305 342 307
rect 344 305 345 307
rect 161 599 162 601
rect 164 599 165 601
rect 161 605 162 607
rect 164 605 165 607
rect 341 19 342 21
rect 344 19 345 21
rect 341 25 342 27
rect 344 25 345 27
rect 301 459 302 461
rect 304 459 305 461
rect 301 465 302 467
rect 304 465 305 467
rect 181 -1 182 1
rect 184 -1 185 1
rect 181 5 182 7
rect 184 5 185 7
rect 101 559 102 561
rect 104 559 105 561
rect 101 565 102 567
rect 104 565 105 567
rect 381 79 382 81
rect 384 79 385 81
rect 381 85 382 87
rect 384 85 385 87
rect 421 -1 422 1
rect 424 -1 425 1
rect 421 5 422 7
rect 424 5 425 7
rect 561 439 562 441
rect 564 439 565 441
rect 561 445 562 447
rect 564 445 565 447
rect 441 479 442 481
rect 444 479 445 481
rect 441 485 442 487
rect 444 485 445 487
rect 301 19 302 21
rect 304 19 305 21
rect 301 25 302 27
rect 304 25 305 27
rect 21 139 22 141
rect 24 139 25 141
rect 21 145 22 147
rect 24 145 25 147
rect 101 39 102 41
rect 104 39 105 41
rect 101 45 102 47
rect 104 45 105 47
rect 521 159 522 161
rect 524 159 525 161
rect 521 165 522 167
rect 524 165 525 167
rect 341 619 342 621
rect 344 619 345 621
rect 341 625 342 627
rect 344 625 345 627
rect 541 259 542 261
rect 544 259 545 261
rect 541 265 542 267
rect 544 265 545 267
rect 421 259 422 261
rect 424 259 425 261
rect 421 265 422 267
rect 424 265 425 267
rect 641 459 642 461
rect 644 459 645 461
rect 641 465 642 467
rect 644 465 645 467
rect 461 319 462 321
rect 464 319 465 321
rect 461 325 462 327
rect 464 325 465 327
rect 301 -1 302 1
rect 304 -1 305 1
rect 301 5 302 7
rect 304 5 305 7
rect 61 319 62 321
rect 64 319 65 321
rect 61 325 62 327
rect 64 325 65 327
rect 301 559 302 561
rect 304 559 305 561
rect 301 565 302 567
rect 304 565 305 567
rect 81 319 82 321
rect 84 319 85 321
rect 81 325 82 327
rect 84 325 85 327
rect 101 199 102 201
rect 104 199 105 201
rect 101 205 102 207
rect 104 205 105 207
rect 161 319 162 321
rect 164 319 165 321
rect 161 325 162 327
rect 164 325 165 327
rect 401 299 402 301
rect 404 299 405 301
rect 401 305 402 307
rect 404 305 405 307
rect 401 479 402 481
rect 404 479 405 481
rect 401 485 402 487
rect 404 485 405 487
rect 61 379 62 381
rect 64 379 65 381
rect 61 385 62 387
rect 64 385 65 387
rect 141 539 142 541
rect 144 539 145 541
rect 141 545 142 547
rect 144 545 145 547
rect 201 599 202 601
rect 204 599 205 601
rect 201 605 202 607
rect 204 605 205 607
rect 221 479 222 481
rect 224 479 225 481
rect 221 485 222 487
rect 224 485 225 487
rect 141 239 142 241
rect 144 239 145 241
rect 141 245 142 247
rect 144 245 145 247
rect 141 19 142 21
rect 144 19 145 21
rect 141 25 142 27
rect 144 25 145 27
rect 201 59 202 61
rect 204 59 205 61
rect 201 65 202 67
rect 204 65 205 67
rect 241 279 242 281
rect 244 279 245 281
rect 241 285 242 287
rect 244 285 245 287
rect 361 239 362 241
rect 364 239 365 241
rect 361 245 362 247
rect 364 245 365 247
rect 481 139 482 141
rect 484 139 485 141
rect 481 145 482 147
rect 484 145 485 147
rect 221 579 222 581
rect 224 579 225 581
rect 221 585 222 587
rect 224 585 225 587
rect 221 459 222 461
rect 224 459 225 461
rect 221 465 222 467
rect 224 465 225 467
rect 241 419 242 421
rect 244 419 245 421
rect 241 425 242 427
rect 244 425 245 427
rect 181 219 182 221
rect 184 219 185 221
rect 181 225 182 227
rect 184 225 185 227
rect 381 619 382 621
rect 384 619 385 621
rect 381 625 382 627
rect 384 625 385 627
rect 1 219 2 221
rect 4 219 5 221
rect 1 225 2 227
rect 4 225 5 227
rect 561 459 562 461
rect 564 459 565 461
rect 561 465 562 467
rect 564 465 565 467
rect 321 339 322 341
rect 324 339 325 341
rect 321 345 322 347
rect 324 345 325 347
rect 41 299 42 301
rect 44 299 45 301
rect 41 305 42 307
rect 44 305 45 307
rect 601 339 602 341
rect 604 339 605 341
rect 601 345 602 347
rect 604 345 605 347
rect 281 599 282 601
rect 284 599 285 601
rect 281 605 282 607
rect 284 605 285 607
rect 581 319 582 321
rect 584 319 585 321
rect 581 325 582 327
rect 584 325 585 327
rect 461 -1 462 1
rect 464 -1 465 1
rect 461 5 462 7
rect 464 5 465 7
rect 241 499 242 501
rect 244 499 245 501
rect 241 505 242 507
rect 244 505 245 507
rect 321 619 322 621
rect 324 619 325 621
rect 321 625 322 627
rect 324 625 325 627
rect 481 519 482 521
rect 484 519 485 521
rect 481 525 482 527
rect 484 525 485 527
rect 401 279 402 281
rect 404 279 405 281
rect 401 285 402 287
rect 404 285 405 287
rect 421 559 422 561
rect 424 559 425 561
rect 421 565 422 567
rect 424 565 425 567
rect 161 399 162 401
rect 164 399 165 401
rect 161 405 162 407
rect 164 405 165 407
rect 401 59 402 61
rect 404 59 405 61
rect 401 65 402 67
rect 404 65 405 67
rect 581 99 582 101
rect 584 99 585 101
rect 581 105 582 107
rect 584 105 585 107
rect 181 299 182 301
rect 184 299 185 301
rect 181 305 182 307
rect 184 305 185 307
rect 1 319 2 321
rect 4 319 5 321
rect 1 325 2 327
rect 4 325 5 327
rect 121 239 122 241
rect 124 239 125 241
rect 121 245 122 247
rect 124 245 125 247
rect 421 19 422 21
rect 424 19 425 21
rect 421 25 422 27
rect 424 25 425 27
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect 161 19 162 21
rect 164 19 165 21
rect 161 25 162 27
rect 164 25 165 27
rect 521 519 522 521
rect 524 519 525 521
rect 521 525 522 527
rect 524 525 525 527
rect 261 599 262 601
rect 264 599 265 601
rect 261 605 262 607
rect 264 605 265 607
rect 561 539 562 541
rect 564 539 565 541
rect 561 545 562 547
rect 564 545 565 547
rect 141 399 142 401
rect 144 399 145 401
rect 141 405 142 407
rect 144 405 145 407
rect 401 619 402 621
rect 404 619 405 621
rect 401 625 402 627
rect 404 625 405 627
rect 641 239 642 241
rect 644 239 645 241
rect 641 245 642 247
rect 644 245 645 247
rect 541 239 542 241
rect 544 239 545 241
rect 541 245 542 247
rect 544 245 545 247
rect 461 479 462 481
rect 464 479 465 481
rect 461 485 462 487
rect 464 485 465 487
rect 21 519 22 521
rect 24 519 25 521
rect 21 525 22 527
rect 24 525 25 527
rect 441 39 442 41
rect 444 39 445 41
rect 441 45 442 47
rect 444 45 445 47
rect 461 359 462 361
rect 464 359 465 361
rect 461 365 462 367
rect 464 365 465 367
rect 61 519 62 521
rect 64 519 65 521
rect 61 525 62 527
rect 64 525 65 527
rect 341 439 342 441
rect 344 439 345 441
rect 341 445 342 447
rect 344 445 345 447
rect 381 119 382 121
rect 384 119 385 121
rect 381 125 382 127
rect 384 125 385 127
rect 81 579 82 581
rect 84 579 85 581
rect 81 585 82 587
rect 84 585 85 587
rect 581 339 582 341
rect 584 339 585 341
rect 581 345 582 347
rect 584 345 585 347
rect 361 219 362 221
rect 364 219 365 221
rect 361 225 362 227
rect 364 225 365 227
rect 441 99 442 101
rect 444 99 445 101
rect 441 105 442 107
rect 444 105 445 107
rect 81 339 82 341
rect 84 339 85 341
rect 81 345 82 347
rect 84 345 85 347
rect 121 19 122 21
rect 124 19 125 21
rect 121 25 122 27
rect 124 25 125 27
rect 301 599 302 601
rect 304 599 305 601
rect 301 605 302 607
rect 304 605 305 607
rect 181 99 182 101
rect 184 99 185 101
rect 181 105 182 107
rect 184 105 185 107
rect 661 199 662 201
rect 664 199 665 201
rect 661 205 662 207
rect 664 205 665 207
rect 21 259 22 261
rect 24 259 25 261
rect 21 265 22 267
rect 24 265 25 267
rect 381 299 382 301
rect 384 299 385 301
rect 381 305 382 307
rect 384 305 385 307
rect 401 239 402 241
rect 404 239 405 241
rect 401 245 402 247
rect 404 245 405 247
rect 61 299 62 301
rect 64 299 65 301
rect 61 305 62 307
rect 64 305 65 307
rect 581 519 582 521
rect 584 519 585 521
rect 581 525 582 527
rect 584 525 585 527
rect 421 619 422 621
rect 424 619 425 621
rect 421 625 422 627
rect 424 625 425 627
rect 21 199 22 201
rect 24 199 25 201
rect 21 205 22 207
rect 24 205 25 207
rect 501 259 502 261
rect 504 259 505 261
rect 501 265 502 267
rect 504 265 505 267
rect 261 219 262 221
rect 264 219 265 221
rect 261 225 262 227
rect 264 225 265 227
rect 81 279 82 281
rect 84 279 85 281
rect 81 285 82 287
rect 84 285 85 287
rect 161 139 162 141
rect 164 139 165 141
rect 161 145 162 147
rect 164 145 165 147
rect 221 419 222 421
rect 224 419 225 421
rect 221 425 222 427
rect 224 425 225 427
rect 121 199 122 201
rect 124 199 125 201
rect 121 205 122 207
rect 124 205 125 207
rect 361 619 362 621
rect 364 619 365 621
rect 361 625 362 627
rect 364 625 365 627
rect 621 259 622 261
rect 624 259 625 261
rect 621 265 622 267
rect 624 265 625 267
rect 61 199 62 201
rect 64 199 65 201
rect 61 205 62 207
rect 64 205 65 207
rect 401 499 402 501
rect 404 499 405 501
rect 401 505 402 507
rect 404 505 405 507
rect 161 -1 162 1
rect 164 -1 165 1
rect 161 5 162 7
rect 164 5 165 7
rect 281 79 282 81
rect 284 79 285 81
rect 281 85 282 87
rect 284 85 285 87
rect 41 179 42 181
rect 44 179 45 181
rect 41 185 42 187
rect 44 185 45 187
rect 661 179 662 181
rect 664 179 665 181
rect 661 185 662 187
rect 664 185 665 187
rect 341 259 342 261
rect 344 259 345 261
rect 341 265 342 267
rect 344 265 345 267
rect 541 359 542 361
rect 544 359 545 361
rect 541 365 542 367
rect 544 365 545 367
rect 81 79 82 81
rect 84 79 85 81
rect 81 85 82 87
rect 84 85 85 87
rect 141 619 142 621
rect 144 619 145 621
rect 141 625 142 627
rect 144 625 145 627
rect 481 79 482 81
rect 484 79 485 81
rect 481 85 482 87
rect 484 85 485 87
rect 161 79 162 81
rect 164 79 165 81
rect 161 85 162 87
rect 164 85 165 87
rect 261 659 262 661
rect 264 659 265 661
rect 261 665 262 667
rect 264 665 265 667
rect 621 439 622 441
rect 624 439 625 441
rect 621 445 622 447
rect 624 445 625 447
rect 101 279 102 281
rect 104 279 105 281
rect 101 285 102 287
rect 104 285 105 287
rect 261 319 262 321
rect 264 319 265 321
rect 261 325 262 327
rect 264 325 265 327
rect 501 399 502 401
rect 504 399 505 401
rect 501 405 502 407
rect 504 405 505 407
rect 181 499 182 501
rect 184 499 185 501
rect 181 505 182 507
rect 184 505 185 507
rect 261 519 262 521
rect 264 519 265 521
rect 261 525 262 527
rect 264 525 265 527
rect 121 459 122 461
rect 124 459 125 461
rect 121 465 122 467
rect 124 465 125 467
rect 621 359 622 361
rect 624 359 625 361
rect 621 365 622 367
rect 624 365 625 367
rect 621 379 622 381
rect 624 379 625 381
rect 621 385 622 387
rect 624 385 625 387
rect 541 179 542 181
rect 544 179 545 181
rect 541 185 542 187
rect 544 185 545 187
rect 181 79 182 81
rect 184 79 185 81
rect 181 85 182 87
rect 184 85 185 87
rect 201 499 202 501
rect 204 499 205 501
rect 201 505 202 507
rect 204 505 205 507
rect 541 99 542 101
rect 544 99 545 101
rect 541 105 542 107
rect 544 105 545 107
rect 261 199 262 201
rect 264 199 265 201
rect 261 205 262 207
rect 264 205 265 207
rect 541 79 542 81
rect 544 79 545 81
rect 541 85 542 87
rect 544 85 545 87
rect 221 339 222 341
rect 224 339 225 341
rect 221 345 222 347
rect 224 345 225 347
rect 581 359 582 361
rect 584 359 585 361
rect 581 365 582 367
rect 584 365 585 367
rect 601 199 602 201
rect 604 199 605 201
rect 601 205 602 207
rect 604 205 605 207
rect 101 159 102 161
rect 104 159 105 161
rect 101 165 102 167
rect 104 165 105 167
rect 41 539 42 541
rect 44 539 45 541
rect 41 545 42 547
rect 44 545 45 547
rect 581 439 582 441
rect 584 439 585 441
rect 581 445 582 447
rect 584 445 585 447
rect 81 519 82 521
rect 84 519 85 521
rect 81 525 82 527
rect 84 525 85 527
rect 141 279 142 281
rect 144 279 145 281
rect 141 285 142 287
rect 144 285 145 287
rect 241 599 242 601
rect 244 599 245 601
rect 241 605 242 607
rect 244 605 245 607
rect 281 259 282 261
rect 284 259 285 261
rect 281 265 282 267
rect 284 265 285 267
rect 161 539 162 541
rect 164 539 165 541
rect 161 545 162 547
rect 164 545 165 547
rect 361 439 362 441
rect 364 439 365 441
rect 361 445 362 447
rect 364 445 365 447
rect 221 79 222 81
rect 224 79 225 81
rect 221 85 222 87
rect 224 85 225 87
rect 401 659 402 661
rect 404 659 405 661
rect 401 665 402 667
rect 404 665 405 667
rect 1 439 2 441
rect 4 439 5 441
rect 1 445 2 447
rect 4 445 5 447
rect 61 459 62 461
rect 64 459 65 461
rect 61 465 62 467
rect 64 465 65 467
rect 541 479 542 481
rect 544 479 545 481
rect 541 485 542 487
rect 544 485 545 487
rect 161 619 162 621
rect 164 619 165 621
rect 161 625 162 627
rect 164 625 165 627
rect 181 579 182 581
rect 184 579 185 581
rect 181 585 182 587
rect 184 585 185 587
rect 1 399 2 401
rect 4 399 5 401
rect 1 405 2 407
rect 4 405 5 407
rect 281 139 282 141
rect 284 139 285 141
rect 281 145 282 147
rect 284 145 285 147
rect 461 279 462 281
rect 464 279 465 281
rect 461 285 462 287
rect 464 285 465 287
rect 421 59 422 61
rect 424 59 425 61
rect 421 65 422 67
rect 424 65 425 67
rect 101 299 102 301
rect 104 299 105 301
rect 101 305 102 307
rect 104 305 105 307
rect 361 119 362 121
rect 364 119 365 121
rect 361 125 362 127
rect 364 125 365 127
rect 1 139 2 141
rect 4 139 5 141
rect 1 145 2 147
rect 4 145 5 147
rect 501 199 502 201
rect 504 199 505 201
rect 501 205 502 207
rect 504 205 505 207
rect 61 259 62 261
rect 64 259 65 261
rect 61 265 62 267
rect 64 265 65 267
rect 401 259 402 261
rect 404 259 405 261
rect 401 265 402 267
rect 404 265 405 267
rect 581 379 582 381
rect 584 379 585 381
rect 581 385 582 387
rect 584 385 585 387
rect 101 599 102 601
rect 104 599 105 601
rect 101 605 102 607
rect 104 605 105 607
rect 601 319 602 321
rect 604 319 605 321
rect 601 325 602 327
rect 604 325 605 327
rect 161 479 162 481
rect 164 479 165 481
rect 161 485 162 487
rect 164 485 165 487
rect 141 419 142 421
rect 144 419 145 421
rect 141 425 142 427
rect 144 425 145 427
rect 261 359 262 361
rect 264 359 265 361
rect 261 365 262 367
rect 264 365 265 367
rect 121 359 122 361
rect 124 359 125 361
rect 121 365 122 367
rect 124 365 125 367
rect 341 279 342 281
rect 344 279 345 281
rect 341 285 342 287
rect 344 285 345 287
rect 101 579 102 581
rect 104 579 105 581
rect 101 585 102 587
rect 104 585 105 587
rect 101 339 102 341
rect 104 339 105 341
rect 101 345 102 347
rect 104 345 105 347
rect 521 459 522 461
rect 524 459 525 461
rect 521 465 522 467
rect 524 465 525 467
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect 621 239 622 241
rect 624 239 625 241
rect 621 245 622 247
rect 624 245 625 247
rect 121 219 122 221
rect 124 219 125 221
rect 121 225 122 227
rect 124 225 125 227
rect 361 19 362 21
rect 364 19 365 21
rect 361 25 362 27
rect 364 25 365 27
rect 381 219 382 221
rect 384 219 385 221
rect 381 225 382 227
rect 384 225 385 227
rect 101 59 102 61
rect 104 59 105 61
rect 101 65 102 67
rect 104 65 105 67
rect 641 399 642 401
rect 644 399 645 401
rect 641 405 642 407
rect 644 405 645 407
rect 41 359 42 361
rect 44 359 45 361
rect 41 365 42 367
rect 44 365 45 367
rect 501 519 502 521
rect 504 519 505 521
rect 501 525 502 527
rect 504 525 505 527
rect 241 159 242 161
rect 244 159 245 161
rect 241 165 242 167
rect 244 165 245 167
rect 621 219 622 221
rect 624 219 625 221
rect 621 225 622 227
rect 624 225 625 227
rect 401 319 402 321
rect 404 319 405 321
rect 401 325 402 327
rect 404 325 405 327
rect 361 59 362 61
rect 364 59 365 61
rect 361 65 362 67
rect 364 65 365 67
rect 601 459 602 461
rect 604 459 605 461
rect 601 465 602 467
rect 604 465 605 467
rect 401 19 402 21
rect 404 19 405 21
rect 401 25 402 27
rect 404 25 405 27
rect 581 219 582 221
rect 584 219 585 221
rect 581 225 582 227
rect 584 225 585 227
rect 481 -1 482 1
rect 484 -1 485 1
rect 481 5 482 7
rect 484 5 485 7
rect 521 119 522 121
rect 524 119 525 121
rect 521 125 522 127
rect 524 125 525 127
rect 601 419 602 421
rect 604 419 605 421
rect 601 425 602 427
rect 604 425 605 427
rect 401 399 402 401
rect 404 399 405 401
rect 401 405 402 407
rect 404 405 405 407
rect 341 39 342 41
rect 344 39 345 41
rect 341 45 342 47
rect 344 45 345 47
rect 321 359 322 361
rect 324 359 325 361
rect 321 365 322 367
rect 324 365 325 367
rect 161 39 162 41
rect 164 39 165 41
rect 161 45 162 47
rect 164 45 165 47
rect 41 159 42 161
rect 44 159 45 161
rect 41 165 42 167
rect 44 165 45 167
rect 121 179 122 181
rect 124 179 125 181
rect 121 185 122 187
rect 124 185 125 187
rect 281 619 282 621
rect 284 619 285 621
rect 281 625 282 627
rect 284 625 285 627
rect 181 599 182 601
rect 184 599 185 601
rect 181 605 182 607
rect 184 605 185 607
rect 581 119 582 121
rect 584 119 585 121
rect 581 125 582 127
rect 584 125 585 127
rect 301 619 302 621
rect 304 619 305 621
rect 301 625 302 627
rect 304 625 305 627
rect 81 379 82 381
rect 84 379 85 381
rect 81 385 82 387
rect 84 385 85 387
rect 641 419 642 421
rect 644 419 645 421
rect 641 425 642 427
rect 644 425 645 427
rect 321 559 322 561
rect 324 559 325 561
rect 321 565 322 567
rect 324 565 325 567
rect 421 339 422 341
rect 424 339 425 341
rect 421 345 422 347
rect 424 345 425 347
rect 61 479 62 481
rect 64 479 65 481
rect 61 485 62 487
rect 64 485 65 487
rect 661 399 662 401
rect 664 399 665 401
rect 661 405 662 407
rect 664 405 665 407
rect 221 19 222 21
rect 224 19 225 21
rect 221 25 222 27
rect 224 25 225 27
rect 1 119 2 121
rect 4 119 5 121
rect 1 125 2 127
rect 4 125 5 127
rect 521 399 522 401
rect 524 399 525 401
rect 521 405 522 407
rect 524 405 525 407
rect 21 479 22 481
rect 24 479 25 481
rect 21 485 22 487
rect 24 485 25 487
rect 181 339 182 341
rect 184 339 185 341
rect 181 345 182 347
rect 184 345 185 347
rect 561 479 562 481
rect 564 479 565 481
rect 561 485 562 487
rect 564 485 565 487
rect 421 179 422 181
rect 424 179 425 181
rect 421 185 422 187
rect 424 185 425 187
rect 281 199 282 201
rect 284 199 285 201
rect 281 205 282 207
rect 284 205 285 207
rect 481 39 482 41
rect 484 39 485 41
rect 481 45 482 47
rect 484 45 485 47
rect 61 219 62 221
rect 64 219 65 221
rect 61 225 62 227
rect 64 225 65 227
rect 141 599 142 601
rect 144 599 145 601
rect 141 605 142 607
rect 144 605 145 607
rect 141 559 142 561
rect 144 559 145 561
rect 141 565 142 567
rect 144 565 145 567
rect 101 119 102 121
rect 104 119 105 121
rect 101 125 102 127
rect 104 125 105 127
rect 481 379 482 381
rect 484 379 485 381
rect 481 385 482 387
rect 484 385 485 387
rect 661 419 662 421
rect 664 419 665 421
rect 661 425 662 427
rect 664 425 665 427
rect 161 59 162 61
rect 164 59 165 61
rect 161 65 162 67
rect 164 65 165 67
rect 1 519 2 521
rect 4 519 5 521
rect 1 525 2 527
rect 4 525 5 527
rect 561 359 562 361
rect 564 359 565 361
rect 561 365 562 367
rect 564 365 565 367
rect 41 119 42 121
rect 44 119 45 121
rect 41 125 42 127
rect 44 125 45 127
rect 141 299 142 301
rect 144 299 145 301
rect 141 305 142 307
rect 144 305 145 307
rect 1 419 2 421
rect 4 419 5 421
rect 1 425 2 427
rect 4 425 5 427
rect 81 219 82 221
rect 84 219 85 221
rect 81 225 82 227
rect 84 225 85 227
rect 21 119 22 121
rect 24 119 25 121
rect 21 125 22 127
rect 24 125 25 127
rect 261 639 262 641
rect 264 639 265 641
rect 261 645 262 647
rect 264 645 265 647
rect 421 479 422 481
rect 424 479 425 481
rect 421 485 422 487
rect 424 485 425 487
rect 381 39 382 41
rect 384 39 385 41
rect 381 45 382 47
rect 384 45 385 47
rect 201 659 202 661
rect 204 659 205 661
rect 201 665 202 667
rect 204 665 205 667
rect 441 499 442 501
rect 444 499 445 501
rect 441 505 442 507
rect 444 505 445 507
rect 461 119 462 121
rect 464 119 465 121
rect 461 125 462 127
rect 464 125 465 127
rect 161 199 162 201
rect 164 199 165 201
rect 161 205 162 207
rect 164 205 165 207
rect 241 39 242 41
rect 244 39 245 41
rect 241 45 242 47
rect 244 45 245 47
rect 301 519 302 521
rect 304 519 305 521
rect 301 525 302 527
rect 304 525 305 527
rect 501 599 502 601
rect 504 599 505 601
rect 501 605 502 607
rect 504 605 505 607
rect 321 259 322 261
rect 324 259 325 261
rect 321 265 322 267
rect 324 265 325 267
rect 601 359 602 361
rect 604 359 605 361
rect 601 365 602 367
rect 604 365 605 367
rect 581 259 582 261
rect 584 259 585 261
rect 581 265 582 267
rect 584 265 585 267
rect 321 659 322 661
rect 324 659 325 661
rect 321 665 322 667
rect 324 665 325 667
rect 561 159 562 161
rect 564 159 565 161
rect 561 165 562 167
rect 564 165 565 167
rect 481 279 482 281
rect 484 279 485 281
rect 481 285 482 287
rect 484 285 485 287
rect 461 539 462 541
rect 464 539 465 541
rect 461 545 462 547
rect 464 545 465 547
rect 1 299 2 301
rect 4 299 5 301
rect 1 305 2 307
rect 4 305 5 307
rect 61 279 62 281
rect 64 279 65 281
rect 61 285 62 287
rect 64 285 65 287
rect 381 319 382 321
rect 384 319 385 321
rect 381 325 382 327
rect 384 325 385 327
rect 121 559 122 561
rect 124 559 125 561
rect 121 565 122 567
rect 124 565 125 567
rect 641 199 642 201
rect 644 199 645 201
rect 641 205 642 207
rect 644 205 645 207
rect 181 419 182 421
rect 184 419 185 421
rect 181 425 182 427
rect 184 425 185 427
rect 381 639 382 641
rect 384 639 385 641
rect 381 645 382 647
rect 384 645 385 647
rect 241 399 242 401
rect 244 399 245 401
rect 241 405 242 407
rect 244 405 245 407
rect 221 399 222 401
rect 224 399 225 401
rect 221 405 222 407
rect 224 405 225 407
rect 201 279 202 281
rect 204 279 205 281
rect 201 285 202 287
rect 204 285 205 287
rect 561 499 562 501
rect 564 499 565 501
rect 561 505 562 507
rect 564 505 565 507
rect 21 419 22 421
rect 24 419 25 421
rect 21 425 22 427
rect 24 425 25 427
rect 461 439 462 441
rect 464 439 465 441
rect 461 445 462 447
rect 464 445 465 447
rect 521 319 522 321
rect 524 319 525 321
rect 521 325 522 327
rect 524 325 525 327
rect 461 299 462 301
rect 464 299 465 301
rect 461 305 462 307
rect 464 305 465 307
rect 281 359 282 361
rect 284 359 285 361
rect 281 365 282 367
rect 284 365 285 367
rect 241 19 242 21
rect 244 19 245 21
rect 241 25 242 27
rect 244 25 245 27
rect 261 279 262 281
rect 264 279 265 281
rect 261 285 262 287
rect 264 285 265 287
rect 241 99 242 101
rect 244 99 245 101
rect 241 105 242 107
rect 244 105 245 107
rect 221 379 222 381
rect 224 379 225 381
rect 221 385 222 387
rect 224 385 225 387
rect 561 239 562 241
rect 564 239 565 241
rect 561 245 562 247
rect 564 245 565 247
rect 521 419 522 421
rect 524 419 525 421
rect 521 425 522 427
rect 524 425 525 427
rect 441 619 442 621
rect 444 619 445 621
rect 441 625 442 627
rect 444 625 445 627
rect 561 339 562 341
rect 564 339 565 341
rect 561 345 562 347
rect 564 345 565 347
rect 181 639 182 641
rect 184 639 185 641
rect 181 645 182 647
rect 184 645 185 647
rect 321 99 322 101
rect 324 99 325 101
rect 321 105 322 107
rect 324 105 325 107
rect 441 279 442 281
rect 444 279 445 281
rect 441 285 442 287
rect 444 285 445 287
rect 621 519 622 521
rect 624 519 625 521
rect 621 525 622 527
rect 624 525 625 527
rect 181 399 182 401
rect 184 399 185 401
rect 181 405 182 407
rect 184 405 185 407
rect 341 559 342 561
rect 344 559 345 561
rect 341 565 342 567
rect 344 565 345 567
rect 301 419 302 421
rect 304 419 305 421
rect 301 425 302 427
rect 304 425 305 427
rect 521 79 522 81
rect 524 79 525 81
rect 521 85 522 87
rect 524 85 525 87
rect 521 499 522 501
rect 524 499 525 501
rect 521 505 522 507
rect 524 505 525 507
rect 101 259 102 261
rect 104 259 105 261
rect 101 265 102 267
rect 104 265 105 267
rect 121 259 122 261
rect 124 259 125 261
rect 121 265 122 267
rect 124 265 125 267
rect 421 199 422 201
rect 424 199 425 201
rect 421 205 422 207
rect 424 205 425 207
rect 141 319 142 321
rect 144 319 145 321
rect 141 325 142 327
rect 144 325 145 327
rect 621 499 622 501
rect 624 499 625 501
rect 621 505 622 507
rect 624 505 625 507
rect 161 339 162 341
rect 164 339 165 341
rect 161 345 162 347
rect 164 345 165 347
rect 201 559 202 561
rect 204 559 205 561
rect 201 565 202 567
rect 204 565 205 567
rect 201 219 202 221
rect 204 219 205 221
rect 201 225 202 227
rect 204 225 205 227
rect 381 499 382 501
rect 384 499 385 501
rect 381 505 382 507
rect 384 505 385 507
rect 521 59 522 61
rect 524 59 525 61
rect 521 65 522 67
rect 524 65 525 67
rect 341 599 342 601
rect 344 599 345 601
rect 341 605 342 607
rect 344 605 345 607
rect 381 159 382 161
rect 384 159 385 161
rect 381 165 382 167
rect 384 165 385 167
rect 161 639 162 641
rect 164 639 165 641
rect 161 645 162 647
rect 164 645 165 647
rect 221 519 222 521
rect 224 519 225 521
rect 221 525 222 527
rect 224 525 225 527
rect 381 419 382 421
rect 384 419 385 421
rect 381 425 382 427
rect 384 425 385 427
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect 501 439 502 441
rect 504 439 505 441
rect 501 445 502 447
rect 504 445 505 447
rect 501 279 502 281
rect 504 279 505 281
rect 501 285 502 287
rect 504 285 505 287
rect 641 339 642 341
rect 644 339 645 341
rect 641 345 642 347
rect 644 345 645 347
rect 141 139 142 141
rect 144 139 145 141
rect 141 145 142 147
rect 144 145 145 147
rect 361 639 362 641
rect 364 639 365 641
rect 361 645 362 647
rect 364 645 365 647
rect 501 479 502 481
rect 504 479 505 481
rect 501 485 502 487
rect 504 485 505 487
rect 381 279 382 281
rect 384 279 385 281
rect 381 285 382 287
rect 384 285 385 287
rect 241 619 242 621
rect 244 619 245 621
rect 241 625 242 627
rect 244 625 245 627
rect 261 559 262 561
rect 264 559 265 561
rect 261 565 262 567
rect 264 565 265 567
rect 101 439 102 441
rect 104 439 105 441
rect 101 445 102 447
rect 104 445 105 447
rect 1 99 2 101
rect 4 99 5 101
rect 1 105 2 107
rect 4 105 5 107
rect 1 199 2 201
rect 4 199 5 201
rect 1 205 2 207
rect 4 205 5 207
rect 261 299 262 301
rect 264 299 265 301
rect 261 305 262 307
rect 264 305 265 307
rect 61 439 62 441
rect 64 439 65 441
rect 61 445 62 447
rect 64 445 65 447
rect 341 -1 342 1
rect 344 -1 345 1
rect 341 5 342 7
rect 344 5 345 7
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect 141 39 142 41
rect 144 39 145 41
rect 141 45 142 47
rect 144 45 145 47
rect 521 259 522 261
rect 524 259 525 261
rect 521 265 522 267
rect 524 265 525 267
rect 441 519 442 521
rect 444 519 445 521
rect 441 525 442 527
rect 444 525 445 527
rect 161 459 162 461
rect 164 459 165 461
rect 161 465 162 467
rect 164 465 165 467
rect 201 519 202 521
rect 204 519 205 521
rect 201 525 202 527
rect 204 525 205 527
rect 541 299 542 301
rect 544 299 545 301
rect 541 305 542 307
rect 544 305 545 307
rect 121 279 122 281
rect 124 279 125 281
rect 121 285 122 287
rect 124 285 125 287
rect 101 319 102 321
rect 104 319 105 321
rect 101 325 102 327
rect 104 325 105 327
rect 421 359 422 361
rect 424 359 425 361
rect 421 365 422 367
rect 424 365 425 367
rect 361 99 362 101
rect 364 99 365 101
rect 361 105 362 107
rect 364 105 365 107
rect 361 339 362 341
rect 364 339 365 341
rect 361 345 362 347
rect 364 345 365 347
rect 321 239 322 241
rect 324 239 325 241
rect 321 245 322 247
rect 324 245 325 247
rect 521 239 522 241
rect 524 239 525 241
rect 521 245 522 247
rect 524 245 525 247
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect 281 479 282 481
rect 284 479 285 481
rect 281 485 282 487
rect 284 485 285 487
rect 601 279 602 281
rect 604 279 605 281
rect 601 285 602 287
rect 604 285 605 287
rect 301 359 302 361
rect 304 359 305 361
rect 301 365 302 367
rect 304 365 305 367
rect 221 139 222 141
rect 224 139 225 141
rect 221 145 222 147
rect 224 145 225 147
rect 201 99 202 101
rect 204 99 205 101
rect 201 105 202 107
rect 204 105 205 107
rect 161 119 162 121
rect 164 119 165 121
rect 161 125 162 127
rect 164 125 165 127
rect 441 379 442 381
rect 444 379 445 381
rect 441 385 442 387
rect 444 385 445 387
rect 121 299 122 301
rect 124 299 125 301
rect 121 305 122 307
rect 124 305 125 307
rect 221 359 222 361
rect 224 359 225 361
rect 221 365 222 367
rect 224 365 225 367
rect 501 579 502 581
rect 504 579 505 581
rect 501 585 502 587
rect 504 585 505 587
rect 501 219 502 221
rect 504 219 505 221
rect 501 225 502 227
rect 504 225 505 227
rect 561 99 562 101
rect 564 99 565 101
rect 561 105 562 107
rect 564 105 565 107
rect 181 439 182 441
rect 184 439 185 441
rect 181 445 182 447
rect 184 445 185 447
rect 1 379 2 381
rect 4 379 5 381
rect 1 385 2 387
rect 4 385 5 387
rect 201 19 202 21
rect 204 19 205 21
rect 201 25 202 27
rect 204 25 205 27
rect 401 159 402 161
rect 404 159 405 161
rect 401 165 402 167
rect 404 165 405 167
rect 461 219 462 221
rect 464 219 465 221
rect 461 225 462 227
rect 464 225 465 227
rect 261 79 262 81
rect 264 79 265 81
rect 261 85 262 87
rect 264 85 265 87
rect 181 619 182 621
rect 184 619 185 621
rect 181 625 182 627
rect 184 625 185 627
rect 361 579 362 581
rect 364 579 365 581
rect 361 585 362 587
rect 364 585 365 587
rect 481 59 482 61
rect 484 59 485 61
rect 481 65 482 67
rect 484 65 485 67
rect 421 139 422 141
rect 424 139 425 141
rect 421 145 422 147
rect 424 145 425 147
rect 561 299 562 301
rect 564 299 565 301
rect 561 305 562 307
rect 564 305 565 307
rect 341 659 342 661
rect 344 659 345 661
rect 341 665 342 667
rect 344 665 345 667
rect 201 139 202 141
rect 204 139 205 141
rect 201 145 202 147
rect 204 145 205 147
rect 561 379 562 381
rect 564 379 565 381
rect 561 385 562 387
rect 564 385 565 387
rect 41 379 42 381
rect 44 379 45 381
rect 41 385 42 387
rect 44 385 45 387
rect 441 19 442 21
rect 444 19 445 21
rect 441 25 442 27
rect 444 25 445 27
rect 601 219 602 221
rect 604 219 605 221
rect 601 225 602 227
rect 604 225 605 227
rect 641 279 642 281
rect 644 279 645 281
rect 641 285 642 287
rect 644 285 645 287
rect 521 379 522 381
rect 524 379 525 381
rect 521 385 522 387
rect 524 385 525 387
rect 201 299 202 301
rect 204 299 205 301
rect 201 305 202 307
rect 204 305 205 307
rect 441 299 442 301
rect 444 299 445 301
rect 441 305 442 307
rect 444 305 445 307
rect 161 99 162 101
rect 164 99 165 101
rect 161 105 162 107
rect 164 105 165 107
rect 101 139 102 141
rect 104 139 105 141
rect 101 145 102 147
rect 104 145 105 147
rect 521 339 522 341
rect 524 339 525 341
rect 521 345 522 347
rect 524 345 525 347
rect 221 -1 222 1
rect 224 -1 225 1
rect 221 5 222 7
rect 224 5 225 7
rect 361 39 362 41
rect 364 39 365 41
rect 361 45 362 47
rect 364 45 365 47
rect 21 319 22 321
rect 24 319 25 321
rect 21 325 22 327
rect 24 325 25 327
rect 41 219 42 221
rect 44 219 45 221
rect 41 225 42 227
rect 44 225 45 227
rect 441 579 442 581
rect 444 579 445 581
rect 441 585 442 587
rect 444 585 445 587
rect 361 139 362 141
rect 364 139 365 141
rect 361 145 362 147
rect 364 145 365 147
rect 401 639 402 641
rect 404 639 405 641
rect 401 645 402 647
rect 404 645 405 647
rect 521 559 522 561
rect 524 559 525 561
rect 521 565 522 567
rect 524 565 525 567
rect 21 339 22 341
rect 24 339 25 341
rect 21 345 22 347
rect 24 345 25 347
rect 541 439 542 441
rect 544 439 545 441
rect 541 445 542 447
rect 544 445 545 447
rect 421 319 422 321
rect 424 319 425 321
rect 421 325 422 327
rect 424 325 425 327
rect 241 79 242 81
rect 244 79 245 81
rect 241 85 242 87
rect 244 85 245 87
rect 561 519 562 521
rect 564 519 565 521
rect 561 525 562 527
rect 564 525 565 527
rect 501 159 502 161
rect 504 159 505 161
rect 501 165 502 167
rect 504 165 505 167
rect 81 419 82 421
rect 84 419 85 421
rect 81 425 82 427
rect 84 425 85 427
rect 201 439 202 441
rect 204 439 205 441
rect 201 445 202 447
rect 204 445 205 447
rect 81 499 82 501
rect 84 499 85 501
rect 81 505 82 507
rect 84 505 85 507
rect 81 539 82 541
rect 84 539 85 541
rect 81 545 82 547
rect 84 545 85 547
rect 61 359 62 361
rect 64 359 65 361
rect 61 365 62 367
rect 64 365 65 367
rect 221 619 222 621
rect 224 619 225 621
rect 221 625 222 627
rect 224 625 225 627
rect 321 419 322 421
rect 324 419 325 421
rect 321 425 322 427
rect 324 425 325 427
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect 161 559 162 561
rect 164 559 165 561
rect 161 565 162 567
rect 164 565 165 567
rect 441 199 442 201
rect 444 199 445 201
rect 441 205 442 207
rect 444 205 445 207
rect 541 319 542 321
rect 544 319 545 321
rect 541 325 542 327
rect 544 325 545 327
rect 621 299 622 301
rect 624 299 625 301
rect 621 305 622 307
rect 624 305 625 307
rect 361 539 362 541
rect 364 539 365 541
rect 361 545 362 547
rect 364 545 365 547
rect 301 659 302 661
rect 304 659 305 661
rect 301 665 302 667
rect 304 665 305 667
rect 441 159 442 161
rect 444 159 445 161
rect 441 165 442 167
rect 444 165 445 167
rect 21 359 22 361
rect 24 359 25 361
rect 21 365 22 367
rect 24 365 25 367
rect 221 219 222 221
rect 224 219 225 221
rect 221 225 222 227
rect 224 225 225 227
rect 161 359 162 361
rect 164 359 165 361
rect 161 365 162 367
rect 164 365 165 367
rect 581 559 582 561
rect 584 559 585 561
rect 581 565 582 567
rect 584 565 585 567
rect 81 239 82 241
rect 84 239 85 241
rect 81 245 82 247
rect 84 245 85 247
rect 201 459 202 461
rect 204 459 205 461
rect 201 465 202 467
rect 204 465 205 467
rect 541 459 542 461
rect 544 459 545 461
rect 541 465 542 467
rect 544 465 545 467
rect 121 519 122 521
rect 124 519 125 521
rect 121 525 122 527
rect 124 525 125 527
rect 501 -1 502 1
rect 504 -1 505 1
rect 501 5 502 7
rect 504 5 505 7
rect 381 379 382 381
rect 384 379 385 381
rect 381 385 382 387
rect 384 385 385 387
rect 481 119 482 121
rect 484 119 485 121
rect 481 125 482 127
rect 484 125 485 127
rect 301 259 302 261
rect 304 259 305 261
rect 301 265 302 267
rect 304 265 305 267
rect 561 279 562 281
rect 564 279 565 281
rect 561 285 562 287
rect 564 285 565 287
rect 341 579 342 581
rect 344 579 345 581
rect 341 585 342 587
rect 344 585 345 587
rect 281 179 282 181
rect 284 179 285 181
rect 281 185 282 187
rect 284 185 285 187
rect 481 219 482 221
rect 484 219 485 221
rect 481 225 482 227
rect 484 225 485 227
rect 181 359 182 361
rect 184 359 185 361
rect 181 365 182 367
rect 184 365 185 367
rect 81 199 82 201
rect 84 199 85 201
rect 81 205 82 207
rect 84 205 85 207
rect 381 239 382 241
rect 384 239 385 241
rect 381 245 382 247
rect 384 245 385 247
rect 1 359 2 361
rect 4 359 5 361
rect 1 365 2 367
rect 4 365 5 367
rect 321 299 322 301
rect 324 299 325 301
rect 321 305 322 307
rect 324 305 325 307
rect 421 519 422 521
rect 424 519 425 521
rect 421 525 422 527
rect 424 525 425 527
rect 381 519 382 521
rect 384 519 385 521
rect 381 525 382 527
rect 384 525 385 527
rect 41 199 42 201
rect 44 199 45 201
rect 41 205 42 207
rect 44 205 45 207
rect 281 39 282 41
rect 284 39 285 41
rect 281 45 282 47
rect 284 45 285 47
rect 281 639 282 641
rect 284 639 285 641
rect 281 645 282 647
rect 284 645 285 647
rect 181 139 182 141
rect 184 139 185 141
rect 181 145 182 147
rect 184 145 185 147
rect 281 279 282 281
rect 284 279 285 281
rect 281 285 282 287
rect 284 285 285 287
rect 321 579 322 581
rect 324 579 325 581
rect 321 585 322 587
rect 324 585 325 587
rect 141 479 142 481
rect 144 479 145 481
rect 141 485 142 487
rect 144 485 145 487
rect 141 459 142 461
rect 144 459 145 461
rect 141 465 142 467
rect 144 465 145 467
rect 61 339 62 341
rect 64 339 65 341
rect 61 345 62 347
rect 64 345 65 347
rect 101 179 102 181
rect 104 179 105 181
rect 101 185 102 187
rect 104 185 105 187
rect 621 479 622 481
rect 624 479 625 481
rect 621 485 622 487
rect 624 485 625 487
rect 401 179 402 181
rect 404 179 405 181
rect 401 185 402 187
rect 404 185 405 187
rect 241 639 242 641
rect 244 639 245 641
rect 241 645 242 647
rect 244 645 245 647
rect 301 239 302 241
rect 304 239 305 241
rect 301 245 302 247
rect 304 245 305 247
rect 321 199 322 201
rect 324 199 325 201
rect 321 205 322 207
rect 324 205 325 207
rect 81 99 82 101
rect 84 99 85 101
rect 81 105 82 107
rect 84 105 85 107
rect 381 199 382 201
rect 384 199 385 201
rect 381 205 382 207
rect 384 205 385 207
rect 501 39 502 41
rect 504 39 505 41
rect 501 45 502 47
rect 504 45 505 47
rect 341 59 342 61
rect 344 59 345 61
rect 341 65 342 67
rect 344 65 345 67
rect 361 359 362 361
rect 364 359 365 361
rect 361 365 362 367
rect 364 365 365 367
rect 581 399 582 401
rect 584 399 585 401
rect 581 405 582 407
rect 584 405 585 407
rect 201 379 202 381
rect 204 379 205 381
rect 201 385 202 387
rect 204 385 205 387
rect 121 599 122 601
rect 124 599 125 601
rect 121 605 122 607
rect 124 605 125 607
rect 41 319 42 321
rect 44 319 45 321
rect 41 325 42 327
rect 44 325 45 327
rect 61 179 62 181
rect 64 179 65 181
rect 61 185 62 187
rect 64 185 65 187
rect 321 599 322 601
rect 324 599 325 601
rect 321 605 322 607
rect 324 605 325 607
rect 101 79 102 81
rect 104 79 105 81
rect 101 85 102 87
rect 104 85 105 87
rect 181 179 182 181
rect 184 179 185 181
rect 181 185 182 187
rect 184 185 185 187
rect 201 419 202 421
rect 204 419 205 421
rect 201 425 202 427
rect 204 425 205 427
rect 421 99 422 101
rect 424 99 425 101
rect 421 105 422 107
rect 424 105 425 107
rect 501 539 502 541
rect 504 539 505 541
rect 501 545 502 547
rect 504 545 505 547
rect 581 419 582 421
rect 584 419 585 421
rect 581 425 582 427
rect 584 425 585 427
rect 561 199 562 201
rect 564 199 565 201
rect 561 205 562 207
rect 564 205 565 207
rect 541 419 542 421
rect 544 419 545 421
rect 541 425 542 427
rect 544 425 545 427
rect 301 319 302 321
rect 304 319 305 321
rect 301 325 302 327
rect 304 325 305 327
rect 261 399 262 401
rect 264 399 265 401
rect 261 405 262 407
rect 264 405 265 407
rect 321 319 322 321
rect 324 319 325 321
rect 321 325 322 327
rect 324 325 325 327
rect 221 539 222 541
rect 224 539 225 541
rect 221 545 222 547
rect 224 545 225 547
rect 421 379 422 381
rect 424 379 425 381
rect 421 385 422 387
rect 424 385 425 387
rect 301 79 302 81
rect 304 79 305 81
rect 301 85 302 87
rect 304 85 305 87
rect 161 379 162 381
rect 164 379 165 381
rect 161 385 162 387
rect 164 385 165 387
rect 161 499 162 501
rect 164 499 165 501
rect 161 505 162 507
rect 164 505 165 507
rect 481 499 482 501
rect 484 499 485 501
rect 481 505 482 507
rect 484 505 485 507
rect 61 79 62 81
rect 64 79 65 81
rect 61 85 62 87
rect 64 85 65 87
rect 481 419 482 421
rect 484 419 485 421
rect 481 425 482 427
rect 484 425 485 427
rect 381 399 382 401
rect 384 399 385 401
rect 381 405 382 407
rect 384 405 385 407
rect 561 139 562 141
rect 564 139 565 141
rect 561 145 562 147
rect 564 145 565 147
rect 201 539 202 541
rect 204 539 205 541
rect 201 545 202 547
rect 204 545 205 547
rect 441 179 442 181
rect 444 179 445 181
rect 441 185 442 187
rect 444 185 445 187
rect 621 419 622 421
rect 624 419 625 421
rect 621 425 622 427
rect 624 425 625 427
rect 181 259 182 261
rect 184 259 185 261
rect 181 265 182 267
rect 184 265 185 267
rect 221 659 222 661
rect 224 659 225 661
rect 221 665 222 667
rect 224 665 225 667
rect 361 419 362 421
rect 364 419 365 421
rect 361 425 362 427
rect 364 425 365 427
rect 121 59 122 61
rect 124 59 125 61
rect 121 65 122 67
rect 124 65 125 67
rect 661 439 662 441
rect 664 439 665 441
rect 661 445 662 447
rect 664 445 665 447
rect 201 339 202 341
rect 204 339 205 341
rect 201 345 202 347
rect 204 345 205 347
rect 541 39 542 41
rect 544 39 545 41
rect 541 45 542 47
rect 544 45 545 47
rect 521 -1 522 1
rect 524 -1 525 1
rect 521 5 522 7
rect 524 5 525 7
rect 581 459 582 461
rect 584 459 585 461
rect 581 465 582 467
rect 584 465 585 467
rect 181 159 182 161
rect 184 159 185 161
rect 181 165 182 167
rect 184 165 185 167
rect 541 119 542 121
rect 544 119 545 121
rect 541 125 542 127
rect 544 125 545 127
rect 421 39 422 41
rect 424 39 425 41
rect 421 45 422 47
rect 424 45 425 47
rect 401 439 402 441
rect 404 439 405 441
rect 401 445 402 447
rect 404 445 405 447
rect 141 359 142 361
rect 144 359 145 361
rect 141 365 142 367
rect 144 365 145 367
rect 441 239 442 241
rect 444 239 445 241
rect 441 245 442 247
rect 444 245 445 247
rect 361 199 362 201
rect 364 199 365 201
rect 361 205 362 207
rect 364 205 365 207
rect 441 559 442 561
rect 444 559 445 561
rect 441 565 442 567
rect 444 565 445 567
rect 181 279 182 281
rect 184 279 185 281
rect 181 285 182 287
rect 184 285 185 287
rect 541 159 542 161
rect 544 159 545 161
rect 541 165 542 167
rect 544 165 545 167
rect 81 359 82 361
rect 84 359 85 361
rect 81 365 82 367
rect 84 365 85 367
rect 241 339 242 341
rect 244 339 245 341
rect 241 345 242 347
rect 244 345 245 347
rect 141 339 142 341
rect 144 339 145 341
rect 141 345 142 347
rect 144 345 145 347
rect 241 559 242 561
rect 244 559 245 561
rect 241 565 242 567
rect 244 565 245 567
rect 301 39 302 41
rect 304 39 305 41
rect 301 45 302 47
rect 304 45 305 47
rect 181 199 182 201
rect 184 199 185 201
rect 181 205 182 207
rect 184 205 185 207
rect 261 459 262 461
rect 264 459 265 461
rect 261 465 262 467
rect 264 465 265 467
rect 421 119 422 121
rect 424 119 425 121
rect 421 125 422 127
rect 424 125 425 127
rect 541 -1 542 1
rect 544 -1 545 1
rect 541 5 542 7
rect 544 5 545 7
rect 281 99 282 101
rect 284 99 285 101
rect 281 105 282 107
rect 284 105 285 107
rect 141 199 142 201
rect 144 199 145 201
rect 141 205 142 207
rect 144 205 145 207
rect 381 -1 382 1
rect 384 -1 385 1
rect 381 5 382 7
rect 384 5 385 7
rect 541 399 542 401
rect 544 399 545 401
rect 541 405 542 407
rect 544 405 545 407
rect 461 39 462 41
rect 464 39 465 41
rect 461 45 462 47
rect 464 45 465 47
rect 381 339 382 341
rect 384 339 385 341
rect 381 345 382 347
rect 384 345 385 347
rect 521 439 522 441
rect 524 439 525 441
rect 521 445 522 447
rect 524 445 525 447
rect 301 99 302 101
rect 304 99 305 101
rect 301 105 302 107
rect 304 105 305 107
rect 241 199 242 201
rect 244 199 245 201
rect 241 205 242 207
rect 244 205 245 207
rect 501 19 502 21
rect 504 19 505 21
rect 501 25 502 27
rect 504 25 505 27
rect 61 539 62 541
rect 64 539 65 541
rect 61 545 62 547
rect 64 545 65 547
rect 161 279 162 281
rect 164 279 165 281
rect 161 285 162 287
rect 164 285 165 287
rect 401 559 402 561
rect 404 559 405 561
rect 401 565 402 567
rect 404 565 405 567
rect 501 319 502 321
rect 504 319 505 321
rect 501 325 502 327
rect 504 325 505 327
rect 121 479 122 481
rect 124 479 125 481
rect 121 485 122 487
rect 124 485 125 487
rect 121 579 122 581
rect 124 579 125 581
rect 121 585 122 587
rect 124 585 125 587
rect 521 599 522 601
rect 524 599 525 601
rect 521 605 522 607
rect 524 605 525 607
rect 541 519 542 521
rect 544 519 545 521
rect 541 525 542 527
rect 544 525 545 527
rect 321 39 322 41
rect 324 39 325 41
rect 321 45 322 47
rect 324 45 325 47
rect 361 559 362 561
rect 364 559 365 561
rect 361 565 362 567
rect 364 565 365 567
rect 301 579 302 581
rect 304 579 305 581
rect 301 585 302 587
rect 304 585 305 587
rect 441 359 442 361
rect 444 359 445 361
rect 441 365 442 367
rect 444 365 445 367
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect 421 299 422 301
rect 424 299 425 301
rect 421 305 422 307
rect 424 305 425 307
rect 361 599 362 601
rect 364 599 365 601
rect 361 605 362 607
rect 364 605 365 607
rect 441 259 442 261
rect 444 259 445 261
rect 441 265 442 267
rect 444 265 445 267
rect 301 159 302 161
rect 304 159 305 161
rect 301 165 302 167
rect 304 165 305 167
rect 221 299 222 301
rect 224 299 225 301
rect 221 305 222 307
rect 224 305 225 307
rect 441 79 442 81
rect 444 79 445 81
rect 441 85 442 87
rect 444 85 445 87
rect 461 619 462 621
rect 464 619 465 621
rect 461 625 462 627
rect 464 625 465 627
rect 201 179 202 181
rect 204 179 205 181
rect 201 185 202 187
rect 204 185 205 187
rect 41 499 42 501
rect 44 499 45 501
rect 41 505 42 507
rect 44 505 45 507
rect 421 539 422 541
rect 424 539 425 541
rect 421 545 422 547
rect 424 545 425 547
rect 141 579 142 581
rect 144 579 145 581
rect 141 585 142 587
rect 144 585 145 587
rect 321 139 322 141
rect 324 139 325 141
rect 321 145 322 147
rect 324 145 325 147
rect 221 199 222 201
rect 224 199 225 201
rect 221 205 222 207
rect 224 205 225 207
rect 121 39 122 41
rect 124 39 125 41
rect 121 45 122 47
rect 124 45 125 47
rect 61 139 62 141
rect 64 139 65 141
rect 61 145 62 147
rect 64 145 65 147
rect 221 639 222 641
rect 224 639 225 641
rect 221 645 222 647
rect 224 645 225 647
rect 601 479 602 481
rect 604 479 605 481
rect 601 485 602 487
rect 604 485 605 487
rect 541 559 542 561
rect 544 559 545 561
rect 541 565 542 567
rect 544 565 545 567
rect 281 219 282 221
rect 284 219 285 221
rect 281 225 282 227
rect 284 225 285 227
rect 1 339 2 341
rect 4 339 5 341
rect 1 345 2 347
rect 4 345 5 347
rect 441 419 442 421
rect 444 419 445 421
rect 441 425 442 427
rect 444 425 445 427
rect 481 299 482 301
rect 484 299 485 301
rect 481 305 482 307
rect 484 305 485 307
rect 1 479 2 481
rect 4 479 5 481
rect 1 485 2 487
rect 4 485 5 487
rect 521 219 522 221
rect 524 219 525 221
rect 521 225 522 227
rect 524 225 525 227
rect 261 19 262 21
rect 264 19 265 21
rect 261 25 262 27
rect 264 25 265 27
rect 461 159 462 161
rect 464 159 465 161
rect 461 165 462 167
rect 464 165 465 167
rect 361 79 362 81
rect 364 79 365 81
rect 361 85 362 87
rect 364 85 365 87
rect 341 419 342 421
rect 344 419 345 421
rect 341 425 342 427
rect 344 425 345 427
rect 301 119 302 121
rect 304 119 305 121
rect 301 125 302 127
rect 304 125 305 127
rect 661 219 662 221
rect 664 219 665 221
rect 661 225 662 227
rect 664 225 665 227
rect 461 599 462 601
rect 464 599 465 601
rect 461 605 462 607
rect 464 605 465 607
rect 581 139 582 141
rect 584 139 585 141
rect 581 145 582 147
rect 584 145 585 147
rect 61 419 62 421
rect 64 419 65 421
rect 61 425 62 427
rect 64 425 65 427
rect 461 99 462 101
rect 464 99 465 101
rect 461 105 462 107
rect 464 105 465 107
rect 561 119 562 121
rect 564 119 565 121
rect 561 125 562 127
rect 564 125 565 127
rect 541 199 542 201
rect 544 199 545 201
rect 541 205 542 207
rect 544 205 545 207
rect 421 499 422 501
rect 424 499 425 501
rect 421 505 422 507
rect 424 505 425 507
rect 301 219 302 221
rect 304 219 305 221
rect 301 225 302 227
rect 304 225 305 227
rect 541 339 542 341
rect 544 339 545 341
rect 541 345 542 347
rect 544 345 545 347
rect 241 439 242 441
rect 244 439 245 441
rect 241 445 242 447
rect 244 445 245 447
rect 481 459 482 461
rect 484 459 485 461
rect 481 465 482 467
rect 484 465 485 467
rect 261 39 262 41
rect 264 39 265 41
rect 261 45 262 47
rect 264 45 265 47
rect 561 419 562 421
rect 564 419 565 421
rect 561 425 562 427
rect 564 425 565 427
rect 341 139 342 141
rect 344 139 345 141
rect 341 145 342 147
rect 344 145 345 147
rect 601 499 602 501
rect 604 499 605 501
rect 601 505 602 507
rect 604 505 605 507
rect 101 419 102 421
rect 104 419 105 421
rect 101 425 102 427
rect 104 425 105 427
rect 521 619 522 621
rect 524 619 525 621
rect 521 625 522 627
rect 524 625 525 627
rect 641 219 642 221
rect 644 219 645 221
rect 641 225 642 227
rect 644 225 645 227
rect 301 59 302 61
rect 304 59 305 61
rect 301 65 302 67
rect 304 65 305 67
rect 241 59 242 61
rect 244 59 245 61
rect 241 65 242 67
rect 244 65 245 67
rect 361 459 362 461
rect 364 459 365 461
rect 361 465 362 467
rect 364 465 365 467
rect 401 599 402 601
rect 404 599 405 601
rect 401 605 402 607
rect 404 605 405 607
rect 501 459 502 461
rect 504 459 505 461
rect 501 465 502 467
rect 504 465 505 467
rect 241 179 242 181
rect 244 179 245 181
rect 241 185 242 187
rect 244 185 245 187
rect 421 579 422 581
rect 424 579 425 581
rect 421 585 422 587
rect 424 585 425 587
rect 201 579 202 581
rect 204 579 205 581
rect 201 585 202 587
rect 204 585 205 587
rect 301 639 302 641
rect 304 639 305 641
rect 301 645 302 647
rect 304 645 305 647
rect 241 359 242 361
rect 244 359 245 361
rect 241 365 242 367
rect 244 365 245 367
rect 501 59 502 61
rect 504 59 505 61
rect 501 65 502 67
rect 504 65 505 67
rect 461 559 462 561
rect 464 559 465 561
rect 461 565 462 567
rect 464 565 465 567
rect 421 239 422 241
rect 424 239 425 241
rect 421 245 422 247
rect 424 245 425 247
rect 341 159 342 161
rect 344 159 345 161
rect 341 165 342 167
rect 344 165 345 167
rect 581 199 582 201
rect 584 199 585 201
rect 581 205 582 207
rect 584 205 585 207
rect 141 219 142 221
rect 144 219 145 221
rect 141 225 142 227
rect 144 225 145 227
rect 341 519 342 521
rect 344 519 345 521
rect 341 525 342 527
rect 344 525 345 527
rect 121 379 122 381
rect 124 379 125 381
rect 121 385 122 387
rect 124 385 125 387
rect 621 319 622 321
rect 624 319 625 321
rect 621 325 622 327
rect 624 325 625 327
rect 121 399 122 401
rect 124 399 125 401
rect 121 405 122 407
rect 124 405 125 407
rect 661 299 662 301
rect 664 299 665 301
rect 661 305 662 307
rect 664 305 665 307
rect 481 199 482 201
rect 484 199 485 201
rect 481 205 482 207
rect 484 205 485 207
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect 141 159 142 161
rect 144 159 145 161
rect 141 165 142 167
rect 144 165 145 167
rect 61 239 62 241
rect 64 239 65 241
rect 61 245 62 247
rect 64 245 65 247
rect 421 459 422 461
rect 424 459 425 461
rect 421 465 422 467
rect 424 465 425 467
rect 221 239 222 241
rect 224 239 225 241
rect 221 245 222 247
rect 224 245 225 247
rect 261 619 262 621
rect 264 619 265 621
rect 261 625 262 627
rect 264 625 265 627
rect 241 239 242 241
rect 244 239 245 241
rect 241 245 242 247
rect 244 245 245 247
rect 81 299 82 301
rect 84 299 85 301
rect 81 305 82 307
rect 84 305 85 307
rect 161 299 162 301
rect 164 299 165 301
rect 161 305 162 307
rect 164 305 165 307
rect 41 519 42 521
rect 44 519 45 521
rect 41 525 42 527
rect 44 525 45 527
rect 521 279 522 281
rect 524 279 525 281
rect 521 285 522 287
rect 524 285 525 287
rect 581 499 582 501
rect 584 499 585 501
rect 581 505 582 507
rect 584 505 585 507
rect 101 379 102 381
rect 104 379 105 381
rect 101 385 102 387
rect 104 385 105 387
rect 221 259 222 261
rect 224 259 225 261
rect 221 265 222 267
rect 224 265 225 267
rect 101 359 102 361
rect 104 359 105 361
rect 101 365 102 367
rect 104 365 105 367
rect 81 139 82 141
rect 84 139 85 141
rect 81 145 82 147
rect 84 145 85 147
rect 41 139 42 141
rect 44 139 45 141
rect 41 145 42 147
rect 44 145 45 147
rect 341 379 342 381
rect 344 379 345 381
rect 341 385 342 387
rect 344 385 345 387
rect 281 499 282 501
rect 284 499 285 501
rect 281 505 282 507
rect 284 505 285 507
rect 641 319 642 321
rect 644 319 645 321
rect 641 325 642 327
rect 644 325 645 327
rect 441 139 442 141
rect 444 139 445 141
rect 441 145 442 147
rect 444 145 445 147
rect 281 159 282 161
rect 284 159 285 161
rect 281 165 282 167
rect 284 165 285 167
rect 141 179 142 181
rect 144 179 145 181
rect 141 185 142 187
rect 144 185 145 187
rect 361 399 362 401
rect 364 399 365 401
rect 361 405 362 407
rect 364 405 365 407
rect 1 179 2 181
rect 4 179 5 181
rect 1 185 2 187
rect 4 185 5 187
rect 481 579 482 581
rect 484 579 485 581
rect 481 585 482 587
rect 484 585 485 587
rect 201 619 202 621
rect 204 619 205 621
rect 201 625 202 627
rect 204 625 205 627
rect 161 579 162 581
rect 164 579 165 581
rect 161 585 162 587
rect 164 585 165 587
rect 181 319 182 321
rect 184 319 185 321
rect 181 325 182 327
rect 184 325 185 327
rect 61 99 62 101
rect 64 99 65 101
rect 61 105 62 107
rect 64 105 65 107
rect 221 119 222 121
rect 224 119 225 121
rect 221 125 222 127
rect 224 125 225 127
<< labels >>
rlabel pdiffusion 423 443 424 444 0 Cellno = 1
rlabel pdiffusion 363 283 364 284 0 Cellno = 2
rlabel pdiffusion 83 483 84 484 0 Cellno = 3
rlabel pdiffusion 123 163 124 164 0 Cellno = 4
rlabel pdiffusion 463 583 464 584 0 Cellno = 5
rlabel pdiffusion 423 163 424 164 0 Cellno = 6
rlabel pdiffusion 523 23 524 24 0 Cellno = 7
rlabel pdiffusion 483 443 484 444 0 Cellno = 8
rlabel pdiffusion 503 183 504 184 0 Cellno = 9
rlabel pdiffusion 383 103 384 104 0 Cellno = 10
rlabel pdiffusion 583 283 584 284 0 Cellno = 11
rlabel pdiffusion 603 243 604 244 0 Cellno = 12
rlabel pdiffusion 323 163 324 164 0 Cellno = 13
rlabel pdiffusion 343 463 344 464 0 Cellno = 14
rlabel pdiffusion 43 283 44 284 0 Cellno = 15
rlabel pdiffusion 263 503 264 504 0 Cellno = 16
rlabel pdiffusion 483 363 484 364 0 Cellno = 17
rlabel pdiffusion 443 323 444 324 0 Cellno = 18
rlabel pdiffusion 283 63 284 64 0 Cellno = 19
rlabel pdiffusion 543 503 544 504 0 Cellno = 20
rlabel pdiffusion 403 363 404 364 0 Cellno = 21
rlabel pdiffusion 463 143 464 144 0 Cellno = 22
rlabel pdiffusion 303 183 304 184 0 Cellno = 23
rlabel pdiffusion 343 243 344 244 0 Cellno = 24
rlabel pdiffusion 203 43 204 44 0 Cellno = 25
rlabel pdiffusion 263 383 264 384 0 Cellno = 26
rlabel pdiffusion 503 563 504 564 0 Cellno = 27
rlabel pdiffusion 223 163 224 164 0 Cellno = 28
rlabel pdiffusion 283 523 284 524 0 Cellno = 29
rlabel pdiffusion 203 483 204 484 0 Cellno = 30
rlabel pdiffusion 463 63 464 64 0 Cellno = 31
rlabel pdiffusion 183 463 184 464 0 Cellno = 32
rlabel pdiffusion 323 23 324 24 0 Cellno = 33
rlabel pdiffusion 323 283 324 284 0 Cellno = 34
rlabel pdiffusion 563 263 564 264 0 Cellno = 35
rlabel pdiffusion 563 323 564 324 0 Cellno = 36
rlabel pdiffusion 663 363 664 364 0 Cellno = 37
rlabel pdiffusion 343 103 344 104 0 Cellno = 38
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 39
rlabel pdiffusion 383 143 384 144 0 Cellno = 40
rlabel pdiffusion 143 383 144 384 0 Cellno = 41
rlabel pdiffusion 323 3 324 4 0 Cellno = 42
rlabel pdiffusion 343 403 344 404 0 Cellno = 43
rlabel pdiffusion 483 403 484 404 0 Cellno = 44
rlabel pdiffusion 163 523 164 524 0 Cellno = 45
rlabel pdiffusion 283 383 284 384 0 Cellno = 46
rlabel pdiffusion 423 423 424 424 0 Cellno = 47
rlabel pdiffusion 543 543 544 544 0 Cellno = 48
rlabel pdiffusion 143 523 144 524 0 Cellno = 49
rlabel pdiffusion 463 203 464 204 0 Cellno = 50
rlabel pdiffusion 383 543 384 544 0 Cellno = 51
rlabel pdiffusion 463 183 464 184 0 Cellno = 52
rlabel pdiffusion 63 403 64 404 0 Cellno = 53
rlabel pdiffusion 243 143 244 144 0 Cellno = 54
rlabel pdiffusion 23 283 24 284 0 Cellno = 55
rlabel pdiffusion 483 603 484 604 0 Cellno = 56
rlabel pdiffusion 383 363 384 364 0 Cellno = 57
rlabel pdiffusion 243 123 244 124 0 Cellno = 58
rlabel pdiffusion 423 643 424 644 0 Cellno = 59
rlabel pdiffusion 603 163 604 164 0 Cellno = 60
rlabel pdiffusion 383 663 384 664 0 Cellno = 61
rlabel pdiffusion 283 123 284 124 0 Cellno = 62
rlabel pdiffusion 303 443 304 444 0 Cellno = 63
rlabel pdiffusion 283 543 284 544 0 Cellno = 64
rlabel pdiffusion 203 83 204 84 0 Cellno = 65
rlabel pdiffusion 23 183 24 184 0 Cellno = 66
rlabel pdiffusion 403 103 404 104 0 Cellno = 67
rlabel pdiffusion 483 643 484 644 0 Cellno = 68
rlabel pdiffusion 363 523 364 524 0 Cellno = 69
rlabel pdiffusion 83 123 84 124 0 Cellno = 70
rlabel pdiffusion 323 123 324 124 0 Cellno = 71
rlabel pdiffusion 303 203 304 204 0 Cellno = 72
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 73
rlabel pdiffusion 303 483 304 484 0 Cellno = 74
rlabel pdiffusion 43 343 44 344 0 Cellno = 75
rlabel pdiffusion 483 243 484 244 0 Cellno = 76
rlabel pdiffusion 203 263 204 264 0 Cellno = 77
rlabel pdiffusion 383 443 384 444 0 Cellno = 78
rlabel pdiffusion 283 303 284 304 0 Cellno = 79
rlabel pdiffusion 623 203 624 204 0 Cellno = 80
rlabel pdiffusion 323 483 324 484 0 Cellno = 81
rlabel pdiffusion 603 523 604 524 0 Cellno = 82
rlabel pdiffusion 123 623 124 624 0 Cellno = 83
rlabel pdiffusion 403 203 404 204 0 Cellno = 84
rlabel pdiffusion 23 403 24 404 0 Cellno = 85
rlabel pdiffusion 283 3 284 4 0 Cellno = 86
rlabel pdiffusion 283 403 284 404 0 Cellno = 87
rlabel pdiffusion 463 243 464 244 0 Cellno = 88
rlabel pdiffusion 303 283 304 284 0 Cellno = 89
rlabel pdiffusion 443 603 444 604 0 Cellno = 90
rlabel pdiffusion 123 423 124 424 0 Cellno = 91
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 92
rlabel pdiffusion 103 543 104 544 0 Cellno = 93
rlabel pdiffusion 343 83 344 84 0 Cellno = 94
rlabel pdiffusion 223 443 224 444 0 Cellno = 95
rlabel pdiffusion 343 183 344 184 0 Cellno = 96
rlabel pdiffusion 363 323 364 324 0 Cellno = 97
rlabel pdiffusion 43 243 44 244 0 Cellno = 98
rlabel pdiffusion 183 663 184 664 0 Cellno = 99
rlabel pdiffusion 523 43 524 44 0 Cellno = 100
rlabel pdiffusion 243 303 244 304 0 Cellno = 101
rlabel pdiffusion 363 163 364 164 0 Cellno = 102
rlabel pdiffusion 403 523 404 524 0 Cellno = 103
rlabel pdiffusion 343 643 344 644 0 Cellno = 104
rlabel pdiffusion 203 163 204 164 0 Cellno = 105
rlabel pdiffusion 23 103 24 104 0 Cellno = 106
rlabel pdiffusion 343 483 344 484 0 Cellno = 107
rlabel pdiffusion 163 263 164 264 0 Cellno = 108
rlabel pdiffusion 503 143 504 144 0 Cellno = 109
rlabel pdiffusion 403 43 404 44 0 Cellno = 110
rlabel pdiffusion 243 543 244 544 0 Cellno = 111
rlabel pdiffusion 523 543 524 544 0 Cellno = 112
rlabel pdiffusion 343 323 344 324 0 Cellno = 113
rlabel pdiffusion 383 463 384 464 0 Cellno = 114
rlabel pdiffusion 103 223 104 224 0 Cellno = 115
rlabel pdiffusion 603 183 604 184 0 Cellno = 116
rlabel pdiffusion 463 343 464 344 0 Cellno = 117
rlabel pdiffusion 83 163 84 164 0 Cellno = 118
rlabel pdiffusion 523 203 524 204 0 Cellno = 119
rlabel pdiffusion 203 363 204 364 0 Cellno = 120
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 121
rlabel pdiffusion 123 143 124 144 0 Cellno = 122
rlabel pdiffusion 163 423 164 424 0 Cellno = 123
rlabel pdiffusion 323 403 324 404 0 Cellno = 124
rlabel pdiffusion 463 523 464 524 0 Cellno = 125
rlabel pdiffusion 363 383 364 384 0 Cellno = 126
rlabel pdiffusion 263 443 264 444 0 Cellno = 127
rlabel pdiffusion 283 443 284 444 0 Cellno = 128
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 129
rlabel pdiffusion 503 383 504 384 0 Cellno = 130
rlabel pdiffusion 503 343 504 344 0 Cellno = 131
rlabel pdiffusion 343 543 344 544 0 Cellno = 132
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 133
rlabel pdiffusion 543 383 544 384 0 Cellno = 134
rlabel pdiffusion 263 263 264 264 0 Cellno = 135
rlabel pdiffusion 443 223 444 224 0 Cellno = 136
rlabel pdiffusion 163 243 164 244 0 Cellno = 137
rlabel pdiffusion 483 543 484 544 0 Cellno = 138
rlabel pdiffusion 383 563 384 564 0 Cellno = 139
rlabel pdiffusion 443 403 444 404 0 Cellno = 140
rlabel pdiffusion 623 183 624 184 0 Cellno = 141
rlabel pdiffusion 303 303 304 304 0 Cellno = 142
rlabel pdiffusion 543 603 544 604 0 Cellno = 143
rlabel pdiffusion 23 243 24 244 0 Cellno = 144
rlabel pdiffusion 323 543 324 544 0 Cellno = 145
rlabel pdiffusion 363 663 364 664 0 Cellno = 146
rlabel pdiffusion 283 343 284 344 0 Cellno = 147
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 148
rlabel pdiffusion 443 463 444 464 0 Cellno = 149
rlabel pdiffusion 263 143 264 144 0 Cellno = 150
rlabel pdiffusion 583 243 584 244 0 Cellno = 151
rlabel pdiffusion 223 63 224 64 0 Cellno = 152
rlabel pdiffusion 403 543 404 544 0 Cellno = 153
rlabel pdiffusion 283 423 284 424 0 Cellno = 154
rlabel pdiffusion 323 503 324 504 0 Cellno = 155
rlabel pdiffusion 323 463 324 464 0 Cellno = 156
rlabel pdiffusion 3 263 4 264 0 Cellno = 157
rlabel pdiffusion 243 463 244 464 0 Cellno = 158
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 159
rlabel pdiffusion 143 123 144 124 0 Cellno = 160
rlabel pdiffusion 563 183 564 184 0 Cellno = 161
rlabel pdiffusion 63 163 64 164 0 Cellno = 162
rlabel pdiffusion 523 143 524 144 0 Cellno = 163
rlabel pdiffusion 263 343 264 344 0 Cellno = 164
rlabel pdiffusion 323 223 324 224 0 Cellno = 165
rlabel pdiffusion 443 443 444 444 0 Cellno = 166
rlabel pdiffusion 203 643 204 644 0 Cellno = 167
rlabel pdiffusion 363 503 364 504 0 Cellno = 168
rlabel pdiffusion 23 503 24 504 0 Cellno = 169
rlabel pdiffusion 383 63 384 64 0 Cellno = 170
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 171
rlabel pdiffusion 343 223 344 224 0 Cellno = 172
rlabel pdiffusion 463 383 464 384 0 Cellno = 173
rlabel pdiffusion 663 283 664 284 0 Cellno = 174
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 175
rlabel pdiffusion 43 263 44 264 0 Cellno = 176
rlabel pdiffusion 243 483 244 484 0 Cellno = 177
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 178
rlabel pdiffusion 663 343 664 344 0 Cellno = 179
rlabel pdiffusion 143 443 144 444 0 Cellno = 180
rlabel pdiffusion 523 103 524 104 0 Cellno = 181
rlabel pdiffusion 623 403 624 404 0 Cellno = 182
rlabel pdiffusion 283 323 284 324 0 Cellno = 183
rlabel pdiffusion 63 123 64 124 0 Cellno = 184
rlabel pdiffusion 343 123 344 124 0 Cellno = 185
rlabel pdiffusion 443 343 444 344 0 Cellno = 186
rlabel pdiffusion 523 363 524 364 0 Cellno = 187
rlabel pdiffusion 323 383 324 384 0 Cellno = 188
rlabel pdiffusion 603 403 604 404 0 Cellno = 189
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 190
rlabel pdiffusion 603 263 604 264 0 Cellno = 191
rlabel pdiffusion 223 43 224 44 0 Cellno = 192
rlabel pdiffusion 123 123 124 124 0 Cellno = 193
rlabel pdiffusion 503 503 504 504 0 Cellno = 194
rlabel pdiffusion 143 503 144 504 0 Cellno = 195
rlabel pdiffusion 443 663 444 664 0 Cellno = 196
rlabel pdiffusion 403 343 404 344 0 Cellno = 197
rlabel pdiffusion 403 223 404 224 0 Cellno = 198
rlabel pdiffusion 123 323 124 324 0 Cellno = 199
rlabel pdiffusion 423 283 424 284 0 Cellno = 200
rlabel pdiffusion 543 223 544 224 0 Cellno = 201
rlabel pdiffusion 223 183 224 184 0 Cellno = 202
rlabel pdiffusion 283 23 284 24 0 Cellno = 203
rlabel pdiffusion 423 603 424 604 0 Cellno = 204
rlabel pdiffusion 183 123 184 124 0 Cellno = 205
rlabel pdiffusion 463 503 464 504 0 Cellno = 206
rlabel pdiffusion 243 383 244 384 0 Cellno = 207
rlabel pdiffusion 243 223 244 224 0 Cellno = 208
rlabel pdiffusion 303 343 304 344 0 Cellno = 209
rlabel pdiffusion 463 263 464 264 0 Cellno = 210
rlabel pdiffusion 123 443 124 444 0 Cellno = 211
rlabel pdiffusion 183 543 184 544 0 Cellno = 212
rlabel pdiffusion 463 83 464 84 0 Cellno = 213
rlabel pdiffusion 583 303 584 304 0 Cellno = 214
rlabel pdiffusion 463 423 464 424 0 Cellno = 215
rlabel pdiffusion 123 343 124 344 0 Cellno = 216
rlabel pdiffusion 223 323 224 324 0 Cellno = 217
rlabel pdiffusion 423 83 424 84 0 Cellno = 218
rlabel pdiffusion 63 563 64 564 0 Cellno = 219
rlabel pdiffusion 423 223 424 224 0 Cellno = 220
rlabel pdiffusion 323 523 324 524 0 Cellno = 221
rlabel pdiffusion 403 143 404 144 0 Cellno = 222
rlabel pdiffusion 403 123 404 124 0 Cellno = 223
rlabel pdiffusion 383 483 384 484 0 Cellno = 224
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 225
rlabel pdiffusion 123 103 124 104 0 Cellno = 226
rlabel pdiffusion 503 103 504 104 0 Cellno = 227
rlabel pdiffusion 303 383 304 384 0 Cellno = 228
rlabel pdiffusion 83 443 84 444 0 Cellno = 229
rlabel pdiffusion 383 603 384 604 0 Cellno = 230
rlabel pdiffusion 203 3 204 4 0 Cellno = 231
rlabel pdiffusion 483 343 484 344 0 Cellno = 232
rlabel pdiffusion 223 103 224 104 0 Cellno = 233
rlabel pdiffusion 163 163 164 164 0 Cellno = 234
rlabel pdiffusion 143 263 144 264 0 Cellno = 235
rlabel pdiffusion 103 503 104 504 0 Cellno = 236
rlabel pdiffusion 163 443 164 444 0 Cellno = 237
rlabel pdiffusion 523 583 524 584 0 Cellno = 238
rlabel pdiffusion 303 543 304 544 0 Cellno = 239
rlabel pdiffusion 383 583 384 584 0 Cellno = 240
rlabel pdiffusion 363 183 364 184 0 Cellno = 241
rlabel pdiffusion 23 223 24 224 0 Cellno = 242
rlabel pdiffusion 663 323 664 324 0 Cellno = 243
rlabel pdiffusion 323 83 324 84 0 Cellno = 244
rlabel pdiffusion 323 63 324 64 0 Cellno = 245
rlabel pdiffusion 263 583 264 584 0 Cellno = 246
rlabel pdiffusion 263 63 264 64 0 Cellno = 247
rlabel pdiffusion 223 503 224 504 0 Cellno = 248
rlabel pdiffusion 463 23 464 24 0 Cellno = 249
rlabel pdiffusion 103 403 104 404 0 Cellno = 250
rlabel pdiffusion 383 23 384 24 0 Cellno = 251
rlabel pdiffusion 263 123 264 124 0 Cellno = 252
rlabel pdiffusion 163 183 164 184 0 Cellno = 253
rlabel pdiffusion 343 203 344 204 0 Cellno = 254
rlabel pdiffusion 503 83 504 84 0 Cellno = 255
rlabel pdiffusion 503 363 504 364 0 Cellno = 256
rlabel pdiffusion 583 183 584 184 0 Cellno = 257
rlabel pdiffusion 363 3 364 4 0 Cellno = 258
rlabel pdiffusion 523 183 524 184 0 Cellno = 259
rlabel pdiffusion 503 123 504 124 0 Cellno = 260
rlabel pdiffusion 603 303 604 304 0 Cellno = 261
rlabel pdiffusion 103 523 104 524 0 Cellno = 262
rlabel pdiffusion 103 243 104 244 0 Cellno = 263
rlabel pdiffusion 83 183 84 184 0 Cellno = 264
rlabel pdiffusion 263 423 264 424 0 Cellno = 265
rlabel pdiffusion 323 643 324 644 0 Cellno = 266
rlabel pdiffusion 223 603 224 604 0 Cellno = 267
rlabel pdiffusion 503 243 504 244 0 Cellno = 268
rlabel pdiffusion 103 463 104 464 0 Cellno = 269
rlabel pdiffusion 403 383 404 384 0 Cellno = 270
rlabel pdiffusion 203 203 204 204 0 Cellno = 271
rlabel pdiffusion 303 403 304 404 0 Cellno = 272
rlabel pdiffusion 83 563 84 564 0 Cellno = 273
rlabel pdiffusion 243 263 244 264 0 Cellno = 274
rlabel pdiffusion 603 143 604 144 0 Cellno = 275
rlabel pdiffusion 183 23 184 24 0 Cellno = 276
rlabel pdiffusion 603 123 604 124 0 Cellno = 277
rlabel pdiffusion 83 463 84 464 0 Cellno = 278
rlabel pdiffusion 543 283 544 284 0 Cellno = 279
rlabel pdiffusion 203 123 204 124 0 Cellno = 280
rlabel pdiffusion 43 483 44 484 0 Cellno = 281
rlabel pdiffusion 123 543 124 544 0 Cellno = 282
rlabel pdiffusion 423 663 424 664 0 Cellno = 283
rlabel pdiffusion 503 423 504 424 0 Cellno = 284
rlabel pdiffusion 23 303 24 304 0 Cellno = 285
rlabel pdiffusion 583 483 584 484 0 Cellno = 286
rlabel pdiffusion 143 83 144 84 0 Cellno = 287
rlabel pdiffusion 323 183 324 184 0 Cellno = 288
rlabel pdiffusion 23 383 24 384 0 Cellno = 289
rlabel pdiffusion 43 423 44 424 0 Cellno = 290
rlabel pdiffusion 643 363 644 364 0 Cellno = 291
rlabel pdiffusion 403 83 404 84 0 Cellno = 292
rlabel pdiffusion 3 243 4 244 0 Cellno = 293
rlabel pdiffusion 183 243 184 244 0 Cellno = 294
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 295
rlabel pdiffusion 283 463 284 464 0 Cellno = 296
rlabel pdiffusion 643 263 644 264 0 Cellno = 297
rlabel pdiffusion 563 223 564 224 0 Cellno = 298
rlabel pdiffusion 443 63 444 64 0 Cellno = 299
rlabel pdiffusion 523 483 524 484 0 Cellno = 300
rlabel pdiffusion 263 103 264 104 0 Cellno = 301
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 302
rlabel pdiffusion 263 483 264 484 0 Cellno = 303
rlabel pdiffusion 183 523 184 524 0 Cellno = 304
rlabel pdiffusion 363 263 364 264 0 Cellno = 305
rlabel pdiffusion 323 443 324 444 0 Cellno = 306
rlabel pdiffusion 363 483 364 484 0 Cellno = 307
rlabel pdiffusion 263 163 264 164 0 Cellno = 308
rlabel pdiffusion 663 243 664 244 0 Cellno = 309
rlabel pdiffusion 203 243 204 244 0 Cellno = 310
rlabel pdiffusion 483 323 484 324 0 Cellno = 311
rlabel pdiffusion 123 503 124 504 0 Cellno = 312
rlabel pdiffusion 43 403 44 404 0 Cellno = 313
rlabel pdiffusion 223 283 224 284 0 Cellno = 314
rlabel pdiffusion 283 663 284 664 0 Cellno = 315
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 316
rlabel pdiffusion 623 343 624 344 0 Cellno = 317
rlabel pdiffusion 483 623 484 624 0 Cellno = 318
rlabel pdiffusion 183 483 184 484 0 Cellno = 319
rlabel pdiffusion 643 303 644 304 0 Cellno = 320
rlabel pdiffusion 103 483 104 484 0 Cellno = 321
rlabel pdiffusion 503 303 504 304 0 Cellno = 322
rlabel pdiffusion 183 563 184 564 0 Cellno = 323
rlabel pdiffusion 363 303 364 304 0 Cellno = 324
rlabel pdiffusion 263 243 264 244 0 Cellno = 325
rlabel pdiffusion 43 463 44 464 0 Cellno = 326
rlabel pdiffusion 403 583 404 584 0 Cellno = 327
rlabel pdiffusion 203 403 204 404 0 Cellno = 328
rlabel pdiffusion 643 483 644 484 0 Cellno = 329
rlabel pdiffusion 103 103 104 104 0 Cellno = 330
rlabel pdiffusion 403 423 404 424 0 Cellno = 331
rlabel pdiffusion 523 303 524 304 0 Cellno = 332
rlabel pdiffusion 243 323 244 324 0 Cellno = 333
rlabel pdiffusion 283 563 284 564 0 Cellno = 334
rlabel pdiffusion 43 443 44 444 0 Cellno = 335
rlabel pdiffusion 3 163 4 164 0 Cellno = 336
rlabel pdiffusion 263 183 264 184 0 Cellno = 337
rlabel pdiffusion 403 463 404 464 0 Cellno = 338
rlabel pdiffusion 603 383 604 384 0 Cellno = 339
rlabel pdiffusion 163 223 164 224 0 Cellno = 340
rlabel pdiffusion 223 563 224 564 0 Cellno = 341
rlabel pdiffusion 483 163 484 164 0 Cellno = 342
rlabel pdiffusion 303 503 304 504 0 Cellno = 343
rlabel pdiffusion 83 403 84 404 0 Cellno = 344
rlabel pdiffusion 343 343 344 344 0 Cellno = 345
rlabel pdiffusion 403 3 404 4 0 Cellno = 346
rlabel pdiffusion 483 183 484 184 0 Cellno = 347
rlabel pdiffusion 423 403 424 404 0 Cellno = 348
rlabel pdiffusion 283 583 284 584 0 Cellno = 349
rlabel pdiffusion 443 123 444 124 0 Cellno = 350
rlabel pdiffusion 183 63 184 64 0 Cellno = 351
rlabel pdiffusion 463 403 464 404 0 Cellno = 352
rlabel pdiffusion 563 403 564 404 0 Cellno = 353
rlabel pdiffusion 543 143 544 144 0 Cellno = 354
rlabel pdiffusion 183 383 184 384 0 Cellno = 355
rlabel pdiffusion 603 443 604 444 0 Cellno = 356
rlabel pdiffusion 483 103 484 104 0 Cellno = 357
rlabel pdiffusion 243 523 244 524 0 Cellno = 358
rlabel pdiffusion 243 583 244 584 0 Cellno = 359
rlabel pdiffusion 383 183 384 184 0 Cellno = 360
rlabel pdiffusion 643 383 644 384 0 Cellno = 361
rlabel pdiffusion 343 503 344 504 0 Cellno = 362
rlabel pdiffusion 63 503 64 504 0 Cellno = 363
rlabel pdiffusion 203 323 204 324 0 Cellno = 364
rlabel pdiffusion 583 163 584 164 0 Cellno = 365
rlabel pdiffusion 123 83 124 84 0 Cellno = 366
rlabel pdiffusion 443 543 444 544 0 Cellno = 367
rlabel pdiffusion 143 63 144 64 0 Cellno = 368
rlabel pdiffusion 3 463 4 464 0 Cellno = 369
rlabel pdiffusion 623 283 624 284 0 Cellno = 370
rlabel pdiffusion 483 563 484 564 0 Cellno = 371
rlabel pdiffusion 23 463 24 464 0 Cellno = 372
rlabel pdiffusion 483 263 484 264 0 Cellno = 373
rlabel pdiffusion 263 543 264 544 0 Cellno = 374
rlabel pdiffusion 263 3 264 4 0 Cellno = 375
rlabel pdiffusion 83 263 84 264 0 Cellno = 376
rlabel pdiffusion 483 483 484 484 0 Cellno = 377
rlabel pdiffusion 283 243 284 244 0 Cellno = 378
rlabel pdiffusion 463 643 464 644 0 Cellno = 379
rlabel pdiffusion 463 463 464 464 0 Cellno = 380
rlabel pdiffusion 343 363 344 364 0 Cellno = 381
rlabel pdiffusion 303 143 304 144 0 Cellno = 382
rlabel pdiffusion 663 263 664 264 0 Cellno = 383
rlabel pdiffusion 383 263 384 264 0 Cellno = 384
rlabel pdiffusion 83 63 84 64 0 Cellno = 385
rlabel pdiffusion 343 303 344 304 0 Cellno = 386
rlabel pdiffusion 163 603 164 604 0 Cellno = 387
rlabel pdiffusion 343 23 344 24 0 Cellno = 388
rlabel pdiffusion 303 463 304 464 0 Cellno = 389
rlabel pdiffusion 183 3 184 4 0 Cellno = 390
rlabel pdiffusion 103 563 104 564 0 Cellno = 391
rlabel pdiffusion 383 83 384 84 0 Cellno = 392
rlabel pdiffusion 423 3 424 4 0 Cellno = 393
rlabel pdiffusion 563 443 564 444 0 Cellno = 394
rlabel pdiffusion 443 483 444 484 0 Cellno = 395
rlabel pdiffusion 303 23 304 24 0 Cellno = 396
rlabel pdiffusion 23 143 24 144 0 Cellno = 397
rlabel pdiffusion 103 43 104 44 0 Cellno = 398
rlabel pdiffusion 523 163 524 164 0 Cellno = 399
rlabel pdiffusion 343 623 344 624 0 Cellno = 400
rlabel pdiffusion 543 263 544 264 0 Cellno = 401
rlabel pdiffusion 423 263 424 264 0 Cellno = 402
rlabel pdiffusion 643 463 644 464 0 Cellno = 403
rlabel pdiffusion 463 323 464 324 0 Cellno = 404
rlabel pdiffusion 303 3 304 4 0 Cellno = 405
rlabel pdiffusion 63 323 64 324 0 Cellno = 406
rlabel pdiffusion 303 563 304 564 0 Cellno = 407
rlabel pdiffusion 83 323 84 324 0 Cellno = 408
rlabel pdiffusion 103 203 104 204 0 Cellno = 409
rlabel pdiffusion 163 323 164 324 0 Cellno = 410
rlabel pdiffusion 403 303 404 304 0 Cellno = 411
rlabel pdiffusion 403 483 404 484 0 Cellno = 412
rlabel pdiffusion 63 383 64 384 0 Cellno = 413
rlabel pdiffusion 143 543 144 544 0 Cellno = 414
rlabel pdiffusion 203 603 204 604 0 Cellno = 415
rlabel pdiffusion 223 483 224 484 0 Cellno = 416
rlabel pdiffusion 143 243 144 244 0 Cellno = 417
rlabel pdiffusion 143 23 144 24 0 Cellno = 418
rlabel pdiffusion 203 63 204 64 0 Cellno = 419
rlabel pdiffusion 243 283 244 284 0 Cellno = 420
rlabel pdiffusion 363 243 364 244 0 Cellno = 421
rlabel pdiffusion 483 143 484 144 0 Cellno = 422
rlabel pdiffusion 223 583 224 584 0 Cellno = 423
rlabel pdiffusion 223 463 224 464 0 Cellno = 424
rlabel pdiffusion 243 423 244 424 0 Cellno = 425
rlabel pdiffusion 183 223 184 224 0 Cellno = 426
rlabel pdiffusion 383 623 384 624 0 Cellno = 427
rlabel pdiffusion 3 223 4 224 0 Cellno = 428
rlabel pdiffusion 563 463 564 464 0 Cellno = 429
rlabel pdiffusion 323 343 324 344 0 Cellno = 430
rlabel pdiffusion 43 303 44 304 0 Cellno = 431
rlabel pdiffusion 603 343 604 344 0 Cellno = 432
rlabel pdiffusion 283 603 284 604 0 Cellno = 433
rlabel pdiffusion 583 323 584 324 0 Cellno = 434
rlabel pdiffusion 463 3 464 4 0 Cellno = 435
rlabel pdiffusion 243 503 244 504 0 Cellno = 436
rlabel pdiffusion 323 623 324 624 0 Cellno = 437
rlabel pdiffusion 483 523 484 524 0 Cellno = 438
rlabel pdiffusion 403 283 404 284 0 Cellno = 439
rlabel pdiffusion 423 563 424 564 0 Cellno = 440
rlabel pdiffusion 163 403 164 404 0 Cellno = 441
rlabel pdiffusion 403 63 404 64 0 Cellno = 442
rlabel pdiffusion 583 103 584 104 0 Cellno = 443
rlabel pdiffusion 183 303 184 304 0 Cellno = 444
rlabel pdiffusion 3 323 4 324 0 Cellno = 445
rlabel pdiffusion 123 243 124 244 0 Cellno = 446
rlabel pdiffusion 423 23 424 24 0 Cellno = 447
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 448
rlabel pdiffusion 163 23 164 24 0 Cellno = 449
rlabel pdiffusion 523 523 524 524 0 Cellno = 450
rlabel pdiffusion 263 603 264 604 0 Cellno = 451
rlabel pdiffusion 563 543 564 544 0 Cellno = 452
rlabel pdiffusion 143 403 144 404 0 Cellno = 453
rlabel pdiffusion 403 623 404 624 0 Cellno = 454
rlabel pdiffusion 643 243 644 244 0 Cellno = 455
rlabel pdiffusion 543 243 544 244 0 Cellno = 456
rlabel pdiffusion 463 483 464 484 0 Cellno = 457
rlabel pdiffusion 23 523 24 524 0 Cellno = 458
rlabel pdiffusion 443 43 444 44 0 Cellno = 459
rlabel pdiffusion 463 363 464 364 0 Cellno = 460
rlabel pdiffusion 63 523 64 524 0 Cellno = 461
rlabel pdiffusion 343 443 344 444 0 Cellno = 462
rlabel pdiffusion 383 123 384 124 0 Cellno = 463
rlabel pdiffusion 83 583 84 584 0 Cellno = 464
rlabel pdiffusion 583 343 584 344 0 Cellno = 465
rlabel pdiffusion 363 223 364 224 0 Cellno = 466
rlabel pdiffusion 443 103 444 104 0 Cellno = 467
rlabel pdiffusion 83 343 84 344 0 Cellno = 468
rlabel pdiffusion 123 23 124 24 0 Cellno = 469
rlabel pdiffusion 303 603 304 604 0 Cellno = 470
rlabel pdiffusion 183 103 184 104 0 Cellno = 471
rlabel pdiffusion 663 203 664 204 0 Cellno = 472
rlabel pdiffusion 23 263 24 264 0 Cellno = 473
rlabel pdiffusion 383 303 384 304 0 Cellno = 474
rlabel pdiffusion 403 243 404 244 0 Cellno = 475
rlabel pdiffusion 63 303 64 304 0 Cellno = 476
rlabel pdiffusion 583 523 584 524 0 Cellno = 477
rlabel pdiffusion 423 623 424 624 0 Cellno = 478
rlabel pdiffusion 23 203 24 204 0 Cellno = 479
rlabel pdiffusion 503 263 504 264 0 Cellno = 480
rlabel pdiffusion 263 223 264 224 0 Cellno = 481
rlabel pdiffusion 83 283 84 284 0 Cellno = 482
rlabel pdiffusion 163 143 164 144 0 Cellno = 483
rlabel pdiffusion 223 423 224 424 0 Cellno = 484
rlabel pdiffusion 123 203 124 204 0 Cellno = 485
rlabel pdiffusion 363 623 364 624 0 Cellno = 486
rlabel pdiffusion 623 263 624 264 0 Cellno = 487
rlabel pdiffusion 63 203 64 204 0 Cellno = 488
rlabel pdiffusion 403 503 404 504 0 Cellno = 489
rlabel pdiffusion 163 3 164 4 0 Cellno = 490
rlabel pdiffusion 283 83 284 84 0 Cellno = 491
rlabel pdiffusion 43 183 44 184 0 Cellno = 492
rlabel pdiffusion 663 183 664 184 0 Cellno = 493
rlabel pdiffusion 343 263 344 264 0 Cellno = 494
rlabel pdiffusion 543 363 544 364 0 Cellno = 495
rlabel pdiffusion 83 83 84 84 0 Cellno = 496
rlabel pdiffusion 143 623 144 624 0 Cellno = 497
rlabel pdiffusion 483 83 484 84 0 Cellno = 498
rlabel pdiffusion 163 83 164 84 0 Cellno = 499
rlabel pdiffusion 263 663 264 664 0 Cellno = 500
rlabel pdiffusion 623 443 624 444 0 Cellno = 501
rlabel pdiffusion 103 283 104 284 0 Cellno = 502
rlabel pdiffusion 263 323 264 324 0 Cellno = 503
rlabel pdiffusion 503 403 504 404 0 Cellno = 504
rlabel pdiffusion 183 503 184 504 0 Cellno = 505
rlabel pdiffusion 263 523 264 524 0 Cellno = 506
rlabel pdiffusion 123 463 124 464 0 Cellno = 507
rlabel pdiffusion 623 363 624 364 0 Cellno = 508
rlabel pdiffusion 623 383 624 384 0 Cellno = 509
rlabel pdiffusion 543 183 544 184 0 Cellno = 510
rlabel pdiffusion 183 83 184 84 0 Cellno = 511
rlabel pdiffusion 203 503 204 504 0 Cellno = 512
rlabel pdiffusion 543 103 544 104 0 Cellno = 513
rlabel pdiffusion 263 203 264 204 0 Cellno = 514
rlabel pdiffusion 543 83 544 84 0 Cellno = 515
rlabel pdiffusion 223 343 224 344 0 Cellno = 516
rlabel pdiffusion 583 363 584 364 0 Cellno = 517
rlabel pdiffusion 603 203 604 204 0 Cellno = 518
rlabel pdiffusion 103 163 104 164 0 Cellno = 519
rlabel pdiffusion 43 543 44 544 0 Cellno = 520
rlabel pdiffusion 583 443 584 444 0 Cellno = 521
rlabel pdiffusion 83 523 84 524 0 Cellno = 522
rlabel pdiffusion 143 283 144 284 0 Cellno = 523
rlabel pdiffusion 243 603 244 604 0 Cellno = 524
rlabel pdiffusion 283 263 284 264 0 Cellno = 525
rlabel pdiffusion 163 543 164 544 0 Cellno = 526
rlabel pdiffusion 363 443 364 444 0 Cellno = 527
rlabel pdiffusion 223 83 224 84 0 Cellno = 528
rlabel pdiffusion 403 663 404 664 0 Cellno = 529
rlabel pdiffusion 3 443 4 444 0 Cellno = 530
rlabel pdiffusion 63 463 64 464 0 Cellno = 531
rlabel pdiffusion 543 483 544 484 0 Cellno = 532
rlabel pdiffusion 163 623 164 624 0 Cellno = 533
rlabel pdiffusion 183 583 184 584 0 Cellno = 534
rlabel pdiffusion 3 403 4 404 0 Cellno = 535
rlabel pdiffusion 283 143 284 144 0 Cellno = 536
rlabel pdiffusion 463 283 464 284 0 Cellno = 537
rlabel pdiffusion 423 63 424 64 0 Cellno = 538
rlabel pdiffusion 103 303 104 304 0 Cellno = 539
rlabel pdiffusion 363 123 364 124 0 Cellno = 540
rlabel pdiffusion 3 143 4 144 0 Cellno = 541
rlabel pdiffusion 503 203 504 204 0 Cellno = 542
rlabel pdiffusion 63 263 64 264 0 Cellno = 543
rlabel pdiffusion 403 263 404 264 0 Cellno = 544
rlabel pdiffusion 583 383 584 384 0 Cellno = 545
rlabel pdiffusion 103 603 104 604 0 Cellno = 546
rlabel pdiffusion 603 323 604 324 0 Cellno = 547
rlabel pdiffusion 163 483 164 484 0 Cellno = 548
rlabel pdiffusion 143 423 144 424 0 Cellno = 549
rlabel pdiffusion 263 363 264 364 0 Cellno = 550
rlabel pdiffusion 123 363 124 364 0 Cellno = 551
rlabel pdiffusion 343 283 344 284 0 Cellno = 552
rlabel pdiffusion 103 583 104 584 0 Cellno = 553
rlabel pdiffusion 103 343 104 344 0 Cellno = 554
rlabel pdiffusion 523 463 524 464 0 Cellno = 555
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 556
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 557
rlabel pdiffusion 623 243 624 244 0 Cellno = 558
rlabel pdiffusion 123 223 124 224 0 Cellno = 559
rlabel pdiffusion 363 23 364 24 0 Cellno = 560
rlabel pdiffusion 383 223 384 224 0 Cellno = 561
rlabel pdiffusion 103 63 104 64 0 Cellno = 562
rlabel pdiffusion 643 403 644 404 0 Cellno = 563
rlabel pdiffusion 43 363 44 364 0 Cellno = 564
rlabel pdiffusion 503 523 504 524 0 Cellno = 565
rlabel pdiffusion 243 163 244 164 0 Cellno = 566
rlabel pdiffusion 623 223 624 224 0 Cellno = 567
rlabel pdiffusion 403 323 404 324 0 Cellno = 568
rlabel pdiffusion 363 63 364 64 0 Cellno = 569
rlabel pdiffusion 603 463 604 464 0 Cellno = 570
rlabel pdiffusion 403 23 404 24 0 Cellno = 571
rlabel pdiffusion 583 223 584 224 0 Cellno = 572
rlabel pdiffusion 483 3 484 4 0 Cellno = 573
rlabel pdiffusion 523 123 524 124 0 Cellno = 574
rlabel pdiffusion 603 423 604 424 0 Cellno = 575
rlabel pdiffusion 403 403 404 404 0 Cellno = 576
rlabel pdiffusion 343 43 344 44 0 Cellno = 577
rlabel pdiffusion 323 363 324 364 0 Cellno = 578
rlabel pdiffusion 163 43 164 44 0 Cellno = 579
rlabel pdiffusion 43 163 44 164 0 Cellno = 580
rlabel pdiffusion 123 183 124 184 0 Cellno = 581
rlabel pdiffusion 283 623 284 624 0 Cellno = 582
rlabel pdiffusion 183 603 184 604 0 Cellno = 583
rlabel pdiffusion 583 123 584 124 0 Cellno = 584
rlabel pdiffusion 303 623 304 624 0 Cellno = 585
rlabel pdiffusion 83 383 84 384 0 Cellno = 586
rlabel pdiffusion 643 423 644 424 0 Cellno = 587
rlabel pdiffusion 323 563 324 564 0 Cellno = 588
rlabel pdiffusion 423 343 424 344 0 Cellno = 589
rlabel pdiffusion 63 483 64 484 0 Cellno = 590
rlabel pdiffusion 663 403 664 404 0 Cellno = 591
rlabel pdiffusion 223 23 224 24 0 Cellno = 592
rlabel pdiffusion 3 123 4 124 0 Cellno = 593
rlabel pdiffusion 523 403 524 404 0 Cellno = 594
rlabel pdiffusion 23 483 24 484 0 Cellno = 595
rlabel pdiffusion 183 343 184 344 0 Cellno = 596
rlabel pdiffusion 563 483 564 484 0 Cellno = 597
rlabel pdiffusion 423 183 424 184 0 Cellno = 598
rlabel pdiffusion 283 203 284 204 0 Cellno = 599
rlabel pdiffusion 483 43 484 44 0 Cellno = 600
rlabel pdiffusion 63 223 64 224 0 Cellno = 601
rlabel pdiffusion 143 603 144 604 0 Cellno = 602
rlabel pdiffusion 143 563 144 564 0 Cellno = 603
rlabel pdiffusion 103 123 104 124 0 Cellno = 604
rlabel pdiffusion 483 383 484 384 0 Cellno = 605
rlabel pdiffusion 663 423 664 424 0 Cellno = 606
rlabel pdiffusion 163 63 164 64 0 Cellno = 607
rlabel pdiffusion 3 523 4 524 0 Cellno = 608
rlabel pdiffusion 563 363 564 364 0 Cellno = 609
rlabel pdiffusion 43 123 44 124 0 Cellno = 610
rlabel pdiffusion 143 303 144 304 0 Cellno = 611
rlabel pdiffusion 3 423 4 424 0 Cellno = 612
rlabel pdiffusion 83 223 84 224 0 Cellno = 613
rlabel pdiffusion 23 123 24 124 0 Cellno = 614
rlabel pdiffusion 263 643 264 644 0 Cellno = 615
rlabel pdiffusion 423 483 424 484 0 Cellno = 616
rlabel pdiffusion 383 43 384 44 0 Cellno = 617
rlabel pdiffusion 203 663 204 664 0 Cellno = 618
rlabel pdiffusion 443 503 444 504 0 Cellno = 619
rlabel pdiffusion 463 123 464 124 0 Cellno = 620
rlabel pdiffusion 163 203 164 204 0 Cellno = 621
rlabel pdiffusion 243 43 244 44 0 Cellno = 622
rlabel pdiffusion 303 523 304 524 0 Cellno = 623
rlabel pdiffusion 503 603 504 604 0 Cellno = 624
rlabel pdiffusion 323 263 324 264 0 Cellno = 625
rlabel pdiffusion 603 363 604 364 0 Cellno = 626
rlabel pdiffusion 583 263 584 264 0 Cellno = 627
rlabel pdiffusion 323 663 324 664 0 Cellno = 628
rlabel pdiffusion 563 163 564 164 0 Cellno = 629
rlabel pdiffusion 483 283 484 284 0 Cellno = 630
rlabel pdiffusion 463 543 464 544 0 Cellno = 631
rlabel pdiffusion 3 303 4 304 0 Cellno = 632
rlabel pdiffusion 63 283 64 284 0 Cellno = 633
rlabel pdiffusion 383 323 384 324 0 Cellno = 634
rlabel pdiffusion 123 563 124 564 0 Cellno = 635
rlabel pdiffusion 643 203 644 204 0 Cellno = 636
rlabel pdiffusion 183 423 184 424 0 Cellno = 637
rlabel pdiffusion 383 643 384 644 0 Cellno = 638
rlabel pdiffusion 243 403 244 404 0 Cellno = 639
rlabel pdiffusion 223 403 224 404 0 Cellno = 640
rlabel pdiffusion 203 283 204 284 0 Cellno = 641
rlabel pdiffusion 563 503 564 504 0 Cellno = 642
rlabel pdiffusion 23 423 24 424 0 Cellno = 643
rlabel pdiffusion 463 443 464 444 0 Cellno = 644
rlabel pdiffusion 523 323 524 324 0 Cellno = 645
rlabel pdiffusion 463 303 464 304 0 Cellno = 646
rlabel pdiffusion 283 363 284 364 0 Cellno = 647
rlabel pdiffusion 243 23 244 24 0 Cellno = 648
rlabel pdiffusion 263 283 264 284 0 Cellno = 649
rlabel pdiffusion 243 103 244 104 0 Cellno = 650
rlabel pdiffusion 223 383 224 384 0 Cellno = 651
rlabel pdiffusion 563 243 564 244 0 Cellno = 652
rlabel pdiffusion 523 423 524 424 0 Cellno = 653
rlabel pdiffusion 443 623 444 624 0 Cellno = 654
rlabel pdiffusion 563 343 564 344 0 Cellno = 655
rlabel pdiffusion 183 643 184 644 0 Cellno = 656
rlabel pdiffusion 323 103 324 104 0 Cellno = 657
rlabel pdiffusion 443 283 444 284 0 Cellno = 658
rlabel pdiffusion 623 523 624 524 0 Cellno = 659
rlabel pdiffusion 183 403 184 404 0 Cellno = 660
rlabel pdiffusion 343 563 344 564 0 Cellno = 661
rlabel pdiffusion 303 423 304 424 0 Cellno = 662
rlabel pdiffusion 523 83 524 84 0 Cellno = 663
rlabel pdiffusion 523 503 524 504 0 Cellno = 664
rlabel pdiffusion 103 263 104 264 0 Cellno = 665
rlabel pdiffusion 123 263 124 264 0 Cellno = 666
rlabel pdiffusion 423 203 424 204 0 Cellno = 667
rlabel pdiffusion 143 323 144 324 0 Cellno = 668
rlabel pdiffusion 623 503 624 504 0 Cellno = 669
rlabel pdiffusion 163 343 164 344 0 Cellno = 670
rlabel pdiffusion 203 563 204 564 0 Cellno = 671
rlabel pdiffusion 203 223 204 224 0 Cellno = 672
rlabel pdiffusion 383 503 384 504 0 Cellno = 673
rlabel pdiffusion 523 63 524 64 0 Cellno = 674
rlabel pdiffusion 343 603 344 604 0 Cellno = 675
rlabel pdiffusion 383 163 384 164 0 Cellno = 676
rlabel pdiffusion 163 643 164 644 0 Cellno = 677
rlabel pdiffusion 223 523 224 524 0 Cellno = 678
rlabel pdiffusion 383 423 384 424 0 Cellno = 679
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 680
rlabel pdiffusion 503 443 504 444 0 Cellno = 681
rlabel pdiffusion 503 283 504 284 0 Cellno = 682
rlabel pdiffusion 643 343 644 344 0 Cellno = 683
rlabel pdiffusion 143 143 144 144 0 Cellno = 684
rlabel pdiffusion 363 643 364 644 0 Cellno = 685
rlabel pdiffusion 503 483 504 484 0 Cellno = 686
rlabel pdiffusion 383 283 384 284 0 Cellno = 687
rlabel pdiffusion 243 623 244 624 0 Cellno = 688
rlabel pdiffusion 263 563 264 564 0 Cellno = 689
rlabel pdiffusion 103 443 104 444 0 Cellno = 690
rlabel pdiffusion 3 103 4 104 0 Cellno = 691
rlabel pdiffusion 3 203 4 204 0 Cellno = 692
rlabel pdiffusion 263 303 264 304 0 Cellno = 693
rlabel pdiffusion 63 443 64 444 0 Cellno = 694
rlabel pdiffusion 343 3 344 4 0 Cellno = 695
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 696
rlabel pdiffusion 143 43 144 44 0 Cellno = 697
rlabel pdiffusion 523 263 524 264 0 Cellno = 698
rlabel pdiffusion 443 523 444 524 0 Cellno = 699
rlabel pdiffusion 163 463 164 464 0 Cellno = 700
rlabel pdiffusion 203 523 204 524 0 Cellno = 701
rlabel pdiffusion 543 303 544 304 0 Cellno = 702
rlabel pdiffusion 123 283 124 284 0 Cellno = 703
rlabel pdiffusion 103 323 104 324 0 Cellno = 704
rlabel pdiffusion 423 363 424 364 0 Cellno = 705
rlabel pdiffusion 363 103 364 104 0 Cellno = 706
rlabel pdiffusion 363 343 364 344 0 Cellno = 707
rlabel pdiffusion 323 243 324 244 0 Cellno = 708
rlabel pdiffusion 523 243 524 244 0 Cellno = 709
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 710
rlabel pdiffusion 283 483 284 484 0 Cellno = 711
rlabel pdiffusion 603 283 604 284 0 Cellno = 712
rlabel pdiffusion 303 363 304 364 0 Cellno = 713
rlabel pdiffusion 223 143 224 144 0 Cellno = 714
rlabel pdiffusion 203 103 204 104 0 Cellno = 715
rlabel pdiffusion 163 123 164 124 0 Cellno = 716
rlabel pdiffusion 443 383 444 384 0 Cellno = 717
rlabel pdiffusion 123 303 124 304 0 Cellno = 718
rlabel pdiffusion 223 363 224 364 0 Cellno = 719
rlabel pdiffusion 503 583 504 584 0 Cellno = 720
rlabel pdiffusion 503 223 504 224 0 Cellno = 721
rlabel pdiffusion 563 103 564 104 0 Cellno = 722
rlabel pdiffusion 183 443 184 444 0 Cellno = 723
rlabel pdiffusion 3 383 4 384 0 Cellno = 724
rlabel pdiffusion 203 23 204 24 0 Cellno = 725
rlabel pdiffusion 403 163 404 164 0 Cellno = 726
rlabel pdiffusion 463 223 464 224 0 Cellno = 727
rlabel pdiffusion 263 83 264 84 0 Cellno = 728
rlabel pdiffusion 183 623 184 624 0 Cellno = 729
rlabel pdiffusion 363 583 364 584 0 Cellno = 730
rlabel pdiffusion 483 63 484 64 0 Cellno = 731
rlabel pdiffusion 423 143 424 144 0 Cellno = 732
rlabel pdiffusion 563 303 564 304 0 Cellno = 733
rlabel pdiffusion 343 663 344 664 0 Cellno = 734
rlabel pdiffusion 203 143 204 144 0 Cellno = 735
rlabel pdiffusion 563 383 564 384 0 Cellno = 736
rlabel pdiffusion 43 383 44 384 0 Cellno = 737
rlabel pdiffusion 443 23 444 24 0 Cellno = 738
rlabel pdiffusion 603 223 604 224 0 Cellno = 739
rlabel pdiffusion 643 283 644 284 0 Cellno = 740
rlabel pdiffusion 523 383 524 384 0 Cellno = 741
rlabel pdiffusion 203 303 204 304 0 Cellno = 742
rlabel pdiffusion 443 303 444 304 0 Cellno = 743
rlabel pdiffusion 163 103 164 104 0 Cellno = 744
rlabel pdiffusion 103 143 104 144 0 Cellno = 745
rlabel pdiffusion 523 343 524 344 0 Cellno = 746
rlabel pdiffusion 223 3 224 4 0 Cellno = 747
rlabel pdiffusion 363 43 364 44 0 Cellno = 748
rlabel pdiffusion 23 323 24 324 0 Cellno = 749
rlabel pdiffusion 43 223 44 224 0 Cellno = 750
rlabel pdiffusion 443 583 444 584 0 Cellno = 751
rlabel pdiffusion 363 143 364 144 0 Cellno = 752
rlabel pdiffusion 403 643 404 644 0 Cellno = 753
rlabel pdiffusion 523 563 524 564 0 Cellno = 754
rlabel pdiffusion 23 343 24 344 0 Cellno = 755
rlabel pdiffusion 543 443 544 444 0 Cellno = 756
rlabel pdiffusion 423 323 424 324 0 Cellno = 757
rlabel pdiffusion 243 83 244 84 0 Cellno = 758
rlabel pdiffusion 563 523 564 524 0 Cellno = 759
rlabel pdiffusion 503 163 504 164 0 Cellno = 760
rlabel pdiffusion 83 423 84 424 0 Cellno = 761
rlabel pdiffusion 203 443 204 444 0 Cellno = 762
rlabel pdiffusion 83 503 84 504 0 Cellno = 763
rlabel pdiffusion 83 543 84 544 0 Cellno = 764
rlabel pdiffusion 63 363 64 364 0 Cellno = 765
rlabel pdiffusion 223 623 224 624 0 Cellno = 766
rlabel pdiffusion 323 423 324 424 0 Cellno = 767
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 768
rlabel pdiffusion 163 563 164 564 0 Cellno = 769
rlabel pdiffusion 443 203 444 204 0 Cellno = 770
rlabel pdiffusion 543 323 544 324 0 Cellno = 771
rlabel pdiffusion 623 303 624 304 0 Cellno = 772
rlabel pdiffusion 363 543 364 544 0 Cellno = 773
rlabel pdiffusion 303 663 304 664 0 Cellno = 774
rlabel pdiffusion 443 163 444 164 0 Cellno = 775
rlabel pdiffusion 23 363 24 364 0 Cellno = 776
rlabel pdiffusion 223 223 224 224 0 Cellno = 777
rlabel pdiffusion 163 363 164 364 0 Cellno = 778
rlabel pdiffusion 583 563 584 564 0 Cellno = 779
rlabel pdiffusion 83 243 84 244 0 Cellno = 780
rlabel pdiffusion 203 463 204 464 0 Cellno = 781
rlabel pdiffusion 543 463 544 464 0 Cellno = 782
rlabel pdiffusion 123 523 124 524 0 Cellno = 783
rlabel pdiffusion 503 3 504 4 0 Cellno = 784
rlabel pdiffusion 383 383 384 384 0 Cellno = 785
rlabel pdiffusion 483 123 484 124 0 Cellno = 786
rlabel pdiffusion 303 263 304 264 0 Cellno = 787
rlabel pdiffusion 563 283 564 284 0 Cellno = 788
rlabel pdiffusion 343 583 344 584 0 Cellno = 789
rlabel pdiffusion 283 183 284 184 0 Cellno = 790
rlabel pdiffusion 483 223 484 224 0 Cellno = 791
rlabel pdiffusion 183 363 184 364 0 Cellno = 792
rlabel pdiffusion 83 203 84 204 0 Cellno = 793
rlabel pdiffusion 383 243 384 244 0 Cellno = 794
rlabel pdiffusion 3 363 4 364 0 Cellno = 795
rlabel pdiffusion 323 303 324 304 0 Cellno = 796
rlabel pdiffusion 423 523 424 524 0 Cellno = 797
rlabel pdiffusion 383 523 384 524 0 Cellno = 798
rlabel pdiffusion 43 203 44 204 0 Cellno = 799
rlabel pdiffusion 283 43 284 44 0 Cellno = 800
rlabel pdiffusion 283 643 284 644 0 Cellno = 801
rlabel pdiffusion 183 143 184 144 0 Cellno = 802
rlabel pdiffusion 283 283 284 284 0 Cellno = 803
rlabel pdiffusion 323 583 324 584 0 Cellno = 804
rlabel pdiffusion 143 483 144 484 0 Cellno = 805
rlabel pdiffusion 143 463 144 464 0 Cellno = 806
rlabel pdiffusion 63 343 64 344 0 Cellno = 807
rlabel pdiffusion 103 183 104 184 0 Cellno = 808
rlabel pdiffusion 623 483 624 484 0 Cellno = 809
rlabel pdiffusion 403 183 404 184 0 Cellno = 810
rlabel pdiffusion 243 643 244 644 0 Cellno = 811
rlabel pdiffusion 303 243 304 244 0 Cellno = 812
rlabel pdiffusion 323 203 324 204 0 Cellno = 813
rlabel pdiffusion 83 103 84 104 0 Cellno = 814
rlabel pdiffusion 383 203 384 204 0 Cellno = 815
rlabel pdiffusion 503 43 504 44 0 Cellno = 816
rlabel pdiffusion 343 63 344 64 0 Cellno = 817
rlabel pdiffusion 363 363 364 364 0 Cellno = 818
rlabel pdiffusion 583 403 584 404 0 Cellno = 819
rlabel pdiffusion 203 383 204 384 0 Cellno = 820
rlabel pdiffusion 123 603 124 604 0 Cellno = 821
rlabel pdiffusion 43 323 44 324 0 Cellno = 822
rlabel pdiffusion 63 183 64 184 0 Cellno = 823
rlabel pdiffusion 323 603 324 604 0 Cellno = 824
rlabel pdiffusion 103 83 104 84 0 Cellno = 825
rlabel pdiffusion 183 183 184 184 0 Cellno = 826
rlabel pdiffusion 203 423 204 424 0 Cellno = 827
rlabel pdiffusion 423 103 424 104 0 Cellno = 828
rlabel pdiffusion 503 543 504 544 0 Cellno = 829
rlabel pdiffusion 583 423 584 424 0 Cellno = 830
rlabel pdiffusion 563 203 564 204 0 Cellno = 831
rlabel pdiffusion 543 423 544 424 0 Cellno = 832
rlabel pdiffusion 303 323 304 324 0 Cellno = 833
rlabel pdiffusion 263 403 264 404 0 Cellno = 834
rlabel pdiffusion 323 323 324 324 0 Cellno = 835
rlabel pdiffusion 223 543 224 544 0 Cellno = 836
rlabel pdiffusion 423 383 424 384 0 Cellno = 837
rlabel pdiffusion 303 83 304 84 0 Cellno = 838
rlabel pdiffusion 163 383 164 384 0 Cellno = 839
rlabel pdiffusion 163 503 164 504 0 Cellno = 840
rlabel pdiffusion 483 503 484 504 0 Cellno = 841
rlabel pdiffusion 63 83 64 84 0 Cellno = 842
rlabel pdiffusion 483 423 484 424 0 Cellno = 843
rlabel pdiffusion 383 403 384 404 0 Cellno = 844
rlabel pdiffusion 563 143 564 144 0 Cellno = 845
rlabel pdiffusion 203 543 204 544 0 Cellno = 846
rlabel pdiffusion 443 183 444 184 0 Cellno = 847
rlabel pdiffusion 623 423 624 424 0 Cellno = 848
rlabel pdiffusion 183 263 184 264 0 Cellno = 849
rlabel pdiffusion 223 663 224 664 0 Cellno = 850
rlabel pdiffusion 363 423 364 424 0 Cellno = 851
rlabel pdiffusion 123 63 124 64 0 Cellno = 852
rlabel pdiffusion 663 443 664 444 0 Cellno = 853
rlabel pdiffusion 203 343 204 344 0 Cellno = 854
rlabel pdiffusion 543 43 544 44 0 Cellno = 855
rlabel pdiffusion 523 3 524 4 0 Cellno = 856
rlabel pdiffusion 583 463 584 464 0 Cellno = 857
rlabel pdiffusion 183 163 184 164 0 Cellno = 858
rlabel pdiffusion 543 123 544 124 0 Cellno = 859
rlabel pdiffusion 423 43 424 44 0 Cellno = 860
rlabel pdiffusion 403 443 404 444 0 Cellno = 861
rlabel pdiffusion 143 363 144 364 0 Cellno = 862
rlabel pdiffusion 443 243 444 244 0 Cellno = 863
rlabel pdiffusion 363 203 364 204 0 Cellno = 864
rlabel pdiffusion 443 563 444 564 0 Cellno = 865
rlabel pdiffusion 183 283 184 284 0 Cellno = 866
rlabel pdiffusion 543 163 544 164 0 Cellno = 867
rlabel pdiffusion 83 363 84 364 0 Cellno = 868
rlabel pdiffusion 243 343 244 344 0 Cellno = 869
rlabel pdiffusion 143 343 144 344 0 Cellno = 870
rlabel pdiffusion 243 563 244 564 0 Cellno = 871
rlabel pdiffusion 303 43 304 44 0 Cellno = 872
rlabel pdiffusion 183 203 184 204 0 Cellno = 873
rlabel pdiffusion 263 463 264 464 0 Cellno = 874
rlabel pdiffusion 423 123 424 124 0 Cellno = 875
rlabel pdiffusion 543 3 544 4 0 Cellno = 876
rlabel pdiffusion 283 103 284 104 0 Cellno = 877
rlabel pdiffusion 143 203 144 204 0 Cellno = 878
rlabel pdiffusion 383 3 384 4 0 Cellno = 879
rlabel pdiffusion 543 403 544 404 0 Cellno = 880
rlabel pdiffusion 463 43 464 44 0 Cellno = 881
rlabel pdiffusion 383 343 384 344 0 Cellno = 882
rlabel pdiffusion 523 443 524 444 0 Cellno = 883
rlabel pdiffusion 303 103 304 104 0 Cellno = 884
rlabel pdiffusion 243 203 244 204 0 Cellno = 885
rlabel pdiffusion 503 23 504 24 0 Cellno = 886
rlabel pdiffusion 63 543 64 544 0 Cellno = 887
rlabel pdiffusion 163 283 164 284 0 Cellno = 888
rlabel pdiffusion 403 563 404 564 0 Cellno = 889
rlabel pdiffusion 503 323 504 324 0 Cellno = 890
rlabel pdiffusion 123 483 124 484 0 Cellno = 891
rlabel pdiffusion 123 583 124 584 0 Cellno = 892
rlabel pdiffusion 523 603 524 604 0 Cellno = 893
rlabel pdiffusion 543 523 544 524 0 Cellno = 894
rlabel pdiffusion 323 43 324 44 0 Cellno = 895
rlabel pdiffusion 363 563 364 564 0 Cellno = 896
rlabel pdiffusion 303 583 304 584 0 Cellno = 897
rlabel pdiffusion 443 363 444 364 0 Cellno = 898
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 899
rlabel pdiffusion 423 303 424 304 0 Cellno = 900
rlabel pdiffusion 363 603 364 604 0 Cellno = 901
rlabel pdiffusion 443 263 444 264 0 Cellno = 902
rlabel pdiffusion 303 163 304 164 0 Cellno = 903
rlabel pdiffusion 223 303 224 304 0 Cellno = 904
rlabel pdiffusion 443 83 444 84 0 Cellno = 905
rlabel pdiffusion 463 623 464 624 0 Cellno = 906
rlabel pdiffusion 203 183 204 184 0 Cellno = 907
rlabel pdiffusion 43 503 44 504 0 Cellno = 908
rlabel pdiffusion 423 543 424 544 0 Cellno = 909
rlabel pdiffusion 143 583 144 584 0 Cellno = 910
rlabel pdiffusion 323 143 324 144 0 Cellno = 911
rlabel pdiffusion 223 203 224 204 0 Cellno = 912
rlabel pdiffusion 123 43 124 44 0 Cellno = 913
rlabel pdiffusion 63 143 64 144 0 Cellno = 914
rlabel pdiffusion 223 643 224 644 0 Cellno = 915
rlabel pdiffusion 603 483 604 484 0 Cellno = 916
rlabel pdiffusion 543 563 544 564 0 Cellno = 917
rlabel pdiffusion 283 223 284 224 0 Cellno = 918
rlabel pdiffusion 3 343 4 344 0 Cellno = 919
rlabel pdiffusion 443 423 444 424 0 Cellno = 920
rlabel pdiffusion 483 303 484 304 0 Cellno = 921
rlabel pdiffusion 3 483 4 484 0 Cellno = 922
rlabel pdiffusion 523 223 524 224 0 Cellno = 923
rlabel pdiffusion 263 23 264 24 0 Cellno = 924
rlabel pdiffusion 463 163 464 164 0 Cellno = 925
rlabel pdiffusion 363 83 364 84 0 Cellno = 926
rlabel pdiffusion 343 423 344 424 0 Cellno = 927
rlabel pdiffusion 303 123 304 124 0 Cellno = 928
rlabel pdiffusion 663 223 664 224 0 Cellno = 929
rlabel pdiffusion 463 603 464 604 0 Cellno = 930
rlabel pdiffusion 583 143 584 144 0 Cellno = 931
rlabel pdiffusion 63 423 64 424 0 Cellno = 932
rlabel pdiffusion 463 103 464 104 0 Cellno = 933
rlabel pdiffusion 563 123 564 124 0 Cellno = 934
rlabel pdiffusion 543 203 544 204 0 Cellno = 935
rlabel pdiffusion 423 503 424 504 0 Cellno = 936
rlabel pdiffusion 303 223 304 224 0 Cellno = 937
rlabel pdiffusion 543 343 544 344 0 Cellno = 938
rlabel pdiffusion 243 443 244 444 0 Cellno = 939
rlabel pdiffusion 483 463 484 464 0 Cellno = 940
rlabel pdiffusion 263 43 264 44 0 Cellno = 941
rlabel pdiffusion 563 423 564 424 0 Cellno = 942
rlabel pdiffusion 343 143 344 144 0 Cellno = 943
rlabel pdiffusion 603 503 604 504 0 Cellno = 944
rlabel pdiffusion 103 423 104 424 0 Cellno = 945
rlabel pdiffusion 523 623 524 624 0 Cellno = 946
rlabel pdiffusion 643 223 644 224 0 Cellno = 947
rlabel pdiffusion 303 63 304 64 0 Cellno = 948
rlabel pdiffusion 243 63 244 64 0 Cellno = 949
rlabel pdiffusion 363 463 364 464 0 Cellno = 950
rlabel pdiffusion 403 603 404 604 0 Cellno = 951
rlabel pdiffusion 503 463 504 464 0 Cellno = 952
rlabel pdiffusion 243 183 244 184 0 Cellno = 953
rlabel pdiffusion 423 583 424 584 0 Cellno = 954
rlabel pdiffusion 203 583 204 584 0 Cellno = 955
rlabel pdiffusion 303 643 304 644 0 Cellno = 956
rlabel pdiffusion 243 363 244 364 0 Cellno = 957
rlabel pdiffusion 503 63 504 64 0 Cellno = 958
rlabel pdiffusion 463 563 464 564 0 Cellno = 959
rlabel pdiffusion 423 243 424 244 0 Cellno = 960
rlabel pdiffusion 343 163 344 164 0 Cellno = 961
rlabel pdiffusion 583 203 584 204 0 Cellno = 962
rlabel pdiffusion 143 223 144 224 0 Cellno = 963
rlabel pdiffusion 343 523 344 524 0 Cellno = 964
rlabel pdiffusion 123 383 124 384 0 Cellno = 965
rlabel pdiffusion 623 323 624 324 0 Cellno = 966
rlabel pdiffusion 123 403 124 404 0 Cellno = 967
rlabel pdiffusion 663 303 664 304 0 Cellno = 968
rlabel pdiffusion 483 203 484 204 0 Cellno = 969
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 970
rlabel pdiffusion 143 163 144 164 0 Cellno = 971
rlabel pdiffusion 63 243 64 244 0 Cellno = 972
rlabel pdiffusion 423 463 424 464 0 Cellno = 973
rlabel pdiffusion 223 243 224 244 0 Cellno = 974
rlabel pdiffusion 263 623 264 624 0 Cellno = 975
rlabel pdiffusion 243 243 244 244 0 Cellno = 976
rlabel pdiffusion 83 303 84 304 0 Cellno = 977
rlabel pdiffusion 163 303 164 304 0 Cellno = 978
rlabel pdiffusion 43 523 44 524 0 Cellno = 979
rlabel pdiffusion 523 283 524 284 0 Cellno = 980
rlabel pdiffusion 583 503 584 504 0 Cellno = 981
rlabel pdiffusion 103 383 104 384 0 Cellno = 982
rlabel pdiffusion 223 263 224 264 0 Cellno = 983
rlabel pdiffusion 103 363 104 364 0 Cellno = 984
rlabel pdiffusion 83 143 84 144 0 Cellno = 985
rlabel pdiffusion 43 143 44 144 0 Cellno = 986
rlabel pdiffusion 343 383 344 384 0 Cellno = 987
rlabel pdiffusion 283 503 284 504 0 Cellno = 988
rlabel pdiffusion 643 323 644 324 0 Cellno = 989
rlabel pdiffusion 443 143 444 144 0 Cellno = 990
rlabel pdiffusion 283 163 284 164 0 Cellno = 991
rlabel pdiffusion 143 183 144 184 0 Cellno = 992
rlabel pdiffusion 363 403 364 404 0 Cellno = 993
rlabel pdiffusion 3 183 4 184 0 Cellno = 994
rlabel pdiffusion 483 583 484 584 0 Cellno = 995
rlabel pdiffusion 203 623 204 624 0 Cellno = 996
rlabel pdiffusion 163 583 164 584 0 Cellno = 997
rlabel pdiffusion 183 323 184 324 0 Cellno = 998
rlabel pdiffusion 63 103 64 104 0 Cellno = 999
rlabel pdiffusion 223 123 224 124 0 Cellno = 1000
<< end >>
