magic
tech scmos
timestamp
<< pdiffusion >>
rect 120 320 121 321
rect 122 320 123 321
rect 123 320 124 321
rect 125 320 126 321
rect 120 321 126 325
rect 120 325 121 326
rect 122 325 123 326
rect 123 325 124 326
rect 125 325 126 326
rect 360 240 361 241
rect 362 240 363 241
rect 363 240 364 241
rect 365 240 366 241
rect 360 241 366 245
rect 360 245 361 246
rect 362 245 363 246
rect 363 245 364 246
rect 365 245 366 246
rect 140 320 141 321
rect 142 320 143 321
rect 143 320 144 321
rect 145 320 146 321
rect 140 321 146 325
rect 140 325 141 326
rect 142 325 143 326
rect 143 325 144 326
rect 145 325 146 326
rect 260 360 261 361
rect 262 360 263 361
rect 263 360 264 361
rect 265 360 266 361
rect 260 361 266 365
rect 260 365 261 366
rect 262 365 263 366
rect 263 365 264 366
rect 265 365 266 366
rect 180 380 181 381
rect 182 380 183 381
rect 183 380 184 381
rect 185 380 186 381
rect 180 381 186 385
rect 180 385 181 386
rect 182 385 183 386
rect 183 385 184 386
rect 185 385 186 386
rect 320 240 321 241
rect 322 240 323 241
rect 323 240 324 241
rect 325 240 326 241
rect 320 241 326 245
rect 320 245 321 246
rect 322 245 323 246
rect 323 245 324 246
rect 325 245 326 246
rect 80 400 81 401
rect 82 400 83 401
rect 83 400 84 401
rect 85 400 86 401
rect 80 401 86 405
rect 80 405 81 406
rect 82 405 83 406
rect 83 405 84 406
rect 85 405 86 406
rect 80 300 81 301
rect 82 300 83 301
rect 83 300 84 301
rect 85 300 86 301
rect 80 301 86 305
rect 80 305 81 306
rect 82 305 83 306
rect 83 305 84 306
rect 85 305 86 306
rect 360 160 361 161
rect 362 160 363 161
rect 363 160 364 161
rect 365 160 366 161
rect 360 161 366 165
rect 360 165 361 166
rect 362 165 363 166
rect 363 165 364 166
rect 365 165 366 166
rect 320 200 321 201
rect 322 200 323 201
rect 323 200 324 201
rect 325 200 326 201
rect 320 201 326 205
rect 320 205 321 206
rect 322 205 323 206
rect 323 205 324 206
rect 325 205 326 206
rect 320 320 321 321
rect 322 320 323 321
rect 323 320 324 321
rect 325 320 326 321
rect 320 321 326 325
rect 320 325 321 326
rect 322 325 323 326
rect 323 325 324 326
rect 325 325 326 326
rect 380 160 381 161
rect 382 160 383 161
rect 383 160 384 161
rect 385 160 386 161
rect 380 161 386 165
rect 380 165 381 166
rect 382 165 383 166
rect 383 165 384 166
rect 385 165 386 166
rect 280 400 281 401
rect 282 400 283 401
rect 283 400 284 401
rect 285 400 286 401
rect 280 401 286 405
rect 280 405 281 406
rect 282 405 283 406
rect 283 405 284 406
rect 285 405 286 406
rect 0 140 1 141
rect 2 140 3 141
rect 3 140 4 141
rect 5 140 6 141
rect 0 141 6 145
rect 0 145 1 146
rect 2 145 3 146
rect 3 145 4 146
rect 5 145 6 146
rect 100 340 101 341
rect 102 340 103 341
rect 103 340 104 341
rect 105 340 106 341
rect 100 341 106 345
rect 100 345 101 346
rect 102 345 103 346
rect 103 345 104 346
rect 105 345 106 346
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect 80 280 81 281
rect 82 280 83 281
rect 83 280 84 281
rect 85 280 86 281
rect 80 281 86 285
rect 80 285 81 286
rect 82 285 83 286
rect 83 285 84 286
rect 85 285 86 286
rect 120 360 121 361
rect 122 360 123 361
rect 123 360 124 361
rect 125 360 126 361
rect 120 361 126 365
rect 120 365 121 366
rect 122 365 123 366
rect 123 365 124 366
rect 125 365 126 366
rect 80 160 81 161
rect 82 160 83 161
rect 83 160 84 161
rect 85 160 86 161
rect 80 161 86 165
rect 80 165 81 166
rect 82 165 83 166
rect 83 165 84 166
rect 85 165 86 166
rect 320 220 321 221
rect 322 220 323 221
rect 323 220 324 221
rect 325 220 326 221
rect 320 221 326 225
rect 320 225 321 226
rect 322 225 323 226
rect 323 225 324 226
rect 325 225 326 226
rect 260 440 261 441
rect 262 440 263 441
rect 263 440 264 441
rect 265 440 266 441
rect 260 441 266 445
rect 260 445 261 446
rect 262 445 263 446
rect 263 445 264 446
rect 265 445 266 446
rect 200 280 201 281
rect 202 280 203 281
rect 203 280 204 281
rect 205 280 206 281
rect 200 281 206 285
rect 200 285 201 286
rect 202 285 203 286
rect 203 285 204 286
rect 205 285 206 286
rect 360 260 361 261
rect 362 260 363 261
rect 363 260 364 261
rect 365 260 366 261
rect 360 261 366 265
rect 360 265 361 266
rect 362 265 363 266
rect 363 265 364 266
rect 365 265 366 266
rect 400 240 401 241
rect 402 240 403 241
rect 403 240 404 241
rect 405 240 406 241
rect 400 241 406 245
rect 400 245 401 246
rect 402 245 403 246
rect 403 245 404 246
rect 405 245 406 246
rect 80 120 81 121
rect 82 120 83 121
rect 83 120 84 121
rect 85 120 86 121
rect 80 121 86 125
rect 80 125 81 126
rect 82 125 83 126
rect 83 125 84 126
rect 85 125 86 126
rect 320 400 321 401
rect 322 400 323 401
rect 323 400 324 401
rect 325 400 326 401
rect 320 401 326 405
rect 320 405 321 406
rect 322 405 323 406
rect 323 405 324 406
rect 325 405 326 406
rect 260 300 261 301
rect 262 300 263 301
rect 263 300 264 301
rect 265 300 266 301
rect 260 301 266 305
rect 260 305 261 306
rect 262 305 263 306
rect 263 305 264 306
rect 265 305 266 306
rect 160 300 161 301
rect 162 300 163 301
rect 163 300 164 301
rect 165 300 166 301
rect 160 301 166 305
rect 160 305 161 306
rect 162 305 163 306
rect 163 305 164 306
rect 165 305 166 306
rect 260 40 261 41
rect 262 40 263 41
rect 263 40 264 41
rect 265 40 266 41
rect 260 41 266 45
rect 260 45 261 46
rect 262 45 263 46
rect 263 45 264 46
rect 265 45 266 46
rect 240 260 241 261
rect 242 260 243 261
rect 243 260 244 261
rect 245 260 246 261
rect 240 261 246 265
rect 240 265 241 266
rect 242 265 243 266
rect 243 265 244 266
rect 245 265 246 266
rect 180 120 181 121
rect 182 120 183 121
rect 183 120 184 121
rect 185 120 186 121
rect 180 121 186 125
rect 180 125 181 126
rect 182 125 183 126
rect 183 125 184 126
rect 185 125 186 126
rect 40 140 41 141
rect 42 140 43 141
rect 43 140 44 141
rect 45 140 46 141
rect 40 141 46 145
rect 40 145 41 146
rect 42 145 43 146
rect 43 145 44 146
rect 45 145 46 146
rect 400 260 401 261
rect 402 260 403 261
rect 403 260 404 261
rect 405 260 406 261
rect 400 261 406 265
rect 400 265 401 266
rect 402 265 403 266
rect 403 265 404 266
rect 405 265 406 266
rect 240 300 241 301
rect 242 300 243 301
rect 243 300 244 301
rect 245 300 246 301
rect 240 301 246 305
rect 240 305 241 306
rect 242 305 243 306
rect 243 305 244 306
rect 245 305 246 306
rect 160 180 161 181
rect 162 180 163 181
rect 163 180 164 181
rect 165 180 166 181
rect 160 181 166 185
rect 160 185 161 186
rect 162 185 163 186
rect 163 185 164 186
rect 165 185 166 186
rect 260 340 261 341
rect 262 340 263 341
rect 263 340 264 341
rect 265 340 266 341
rect 260 341 266 345
rect 260 345 261 346
rect 262 345 263 346
rect 263 345 264 346
rect 265 345 266 346
rect 120 240 121 241
rect 122 240 123 241
rect 123 240 124 241
rect 125 240 126 241
rect 120 241 126 245
rect 120 245 121 246
rect 122 245 123 246
rect 123 245 124 246
rect 125 245 126 246
rect 400 160 401 161
rect 402 160 403 161
rect 403 160 404 161
rect 405 160 406 161
rect 400 161 406 165
rect 400 165 401 166
rect 402 165 403 166
rect 403 165 404 166
rect 405 165 406 166
rect 40 160 41 161
rect 42 160 43 161
rect 43 160 44 161
rect 45 160 46 161
rect 40 161 46 165
rect 40 165 41 166
rect 42 165 43 166
rect 43 165 44 166
rect 45 165 46 166
rect 280 380 281 381
rect 282 380 283 381
rect 283 380 284 381
rect 285 380 286 381
rect 280 381 286 385
rect 280 385 281 386
rect 282 385 283 386
rect 283 385 284 386
rect 285 385 286 386
rect 140 400 141 401
rect 142 400 143 401
rect 143 400 144 401
rect 145 400 146 401
rect 140 401 146 405
rect 140 405 141 406
rect 142 405 143 406
rect 143 405 144 406
rect 145 405 146 406
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect 280 100 281 101
rect 282 100 283 101
rect 283 100 284 101
rect 285 100 286 101
rect 280 101 286 105
rect 280 105 281 106
rect 282 105 283 106
rect 283 105 284 106
rect 285 105 286 106
rect 100 80 101 81
rect 102 80 103 81
rect 103 80 104 81
rect 105 80 106 81
rect 100 81 106 85
rect 100 85 101 86
rect 102 85 103 86
rect 103 85 104 86
rect 105 85 106 86
rect 400 200 401 201
rect 402 200 403 201
rect 403 200 404 201
rect 405 200 406 201
rect 400 201 406 205
rect 400 205 401 206
rect 402 205 403 206
rect 403 205 404 206
rect 405 205 406 206
rect 280 300 281 301
rect 282 300 283 301
rect 283 300 284 301
rect 285 300 286 301
rect 280 301 286 305
rect 280 305 281 306
rect 282 305 283 306
rect 283 305 284 306
rect 285 305 286 306
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect 280 440 281 441
rect 282 440 283 441
rect 283 440 284 441
rect 285 440 286 441
rect 280 441 286 445
rect 280 445 281 446
rect 282 445 283 446
rect 283 445 284 446
rect 285 445 286 446
rect 160 340 161 341
rect 162 340 163 341
rect 163 340 164 341
rect 165 340 166 341
rect 160 341 166 345
rect 160 345 161 346
rect 162 345 163 346
rect 163 345 164 346
rect 165 345 166 346
rect 100 100 101 101
rect 102 100 103 101
rect 103 100 104 101
rect 105 100 106 101
rect 100 101 106 105
rect 100 105 101 106
rect 102 105 103 106
rect 103 105 104 106
rect 105 105 106 106
rect 200 220 201 221
rect 202 220 203 221
rect 203 220 204 221
rect 205 220 206 221
rect 200 221 206 225
rect 200 225 201 226
rect 202 225 203 226
rect 203 225 204 226
rect 205 225 206 226
rect 100 320 101 321
rect 102 320 103 321
rect 103 320 104 321
rect 105 320 106 321
rect 100 321 106 325
rect 100 325 101 326
rect 102 325 103 326
rect 103 325 104 326
rect 105 325 106 326
rect 160 260 161 261
rect 162 260 163 261
rect 163 260 164 261
rect 165 260 166 261
rect 160 261 166 265
rect 160 265 161 266
rect 162 265 163 266
rect 163 265 164 266
rect 165 265 166 266
rect 120 200 121 201
rect 122 200 123 201
rect 123 200 124 201
rect 125 200 126 201
rect 120 201 126 205
rect 120 205 121 206
rect 122 205 123 206
rect 123 205 124 206
rect 125 205 126 206
rect 280 60 281 61
rect 282 60 283 61
rect 283 60 284 61
rect 285 60 286 61
rect 280 61 286 65
rect 280 65 281 66
rect 282 65 283 66
rect 283 65 284 66
rect 285 65 286 66
rect 80 320 81 321
rect 82 320 83 321
rect 83 320 84 321
rect 85 320 86 321
rect 80 321 86 325
rect 80 325 81 326
rect 82 325 83 326
rect 83 325 84 326
rect 85 325 86 326
rect 360 360 361 361
rect 362 360 363 361
rect 363 360 364 361
rect 365 360 366 361
rect 360 361 366 365
rect 360 365 361 366
rect 362 365 363 366
rect 363 365 364 366
rect 365 365 366 366
rect 200 120 201 121
rect 202 120 203 121
rect 203 120 204 121
rect 205 120 206 121
rect 200 121 206 125
rect 200 125 201 126
rect 202 125 203 126
rect 203 125 204 126
rect 205 125 206 126
rect 240 280 241 281
rect 242 280 243 281
rect 243 280 244 281
rect 245 280 246 281
rect 240 281 246 285
rect 240 285 241 286
rect 242 285 243 286
rect 243 285 244 286
rect 245 285 246 286
rect 260 220 261 221
rect 262 220 263 221
rect 263 220 264 221
rect 265 220 266 221
rect 260 221 266 225
rect 260 225 261 226
rect 262 225 263 226
rect 263 225 264 226
rect 265 225 266 226
rect 220 200 221 201
rect 222 200 223 201
rect 223 200 224 201
rect 225 200 226 201
rect 220 201 226 205
rect 220 205 221 206
rect 222 205 223 206
rect 223 205 224 206
rect 225 205 226 206
rect 260 400 261 401
rect 262 400 263 401
rect 263 400 264 401
rect 265 400 266 401
rect 260 401 266 405
rect 260 405 261 406
rect 262 405 263 406
rect 263 405 264 406
rect 265 405 266 406
rect 140 240 141 241
rect 142 240 143 241
rect 143 240 144 241
rect 145 240 146 241
rect 140 241 146 245
rect 140 245 141 246
rect 142 245 143 246
rect 143 245 144 246
rect 145 245 146 246
rect 240 160 241 161
rect 242 160 243 161
rect 243 160 244 161
rect 245 160 246 161
rect 240 161 246 165
rect 240 165 241 166
rect 242 165 243 166
rect 243 165 244 166
rect 245 165 246 166
rect 100 240 101 241
rect 102 240 103 241
rect 103 240 104 241
rect 105 240 106 241
rect 100 241 106 245
rect 100 245 101 246
rect 102 245 103 246
rect 103 245 104 246
rect 105 245 106 246
rect 160 320 161 321
rect 162 320 163 321
rect 163 320 164 321
rect 165 320 166 321
rect 160 321 166 325
rect 160 325 161 326
rect 162 325 163 326
rect 163 325 164 326
rect 165 325 166 326
rect 160 160 161 161
rect 162 160 163 161
rect 163 160 164 161
rect 165 160 166 161
rect 160 161 166 165
rect 160 165 161 166
rect 162 165 163 166
rect 163 165 164 166
rect 165 165 166 166
rect 80 360 81 361
rect 82 360 83 361
rect 83 360 84 361
rect 85 360 86 361
rect 80 361 86 365
rect 80 365 81 366
rect 82 365 83 366
rect 83 365 84 366
rect 85 365 86 366
rect 40 100 41 101
rect 42 100 43 101
rect 43 100 44 101
rect 45 100 46 101
rect 40 101 46 105
rect 40 105 41 106
rect 42 105 43 106
rect 43 105 44 106
rect 45 105 46 106
rect 200 440 201 441
rect 202 440 203 441
rect 203 440 204 441
rect 205 440 206 441
rect 200 441 206 445
rect 200 445 201 446
rect 202 445 203 446
rect 203 445 204 446
rect 205 445 206 446
rect 60 200 61 201
rect 62 200 63 201
rect 63 200 64 201
rect 65 200 66 201
rect 60 201 66 205
rect 60 205 61 206
rect 62 205 63 206
rect 63 205 64 206
rect 65 205 66 206
rect 0 180 1 181
rect 2 180 3 181
rect 3 180 4 181
rect 5 180 6 181
rect 0 181 6 185
rect 0 185 1 186
rect 2 185 3 186
rect 3 185 4 186
rect 5 185 6 186
rect 180 200 181 201
rect 182 200 183 201
rect 183 200 184 201
rect 185 200 186 201
rect 180 201 186 205
rect 180 205 181 206
rect 182 205 183 206
rect 183 205 184 206
rect 185 205 186 206
rect 300 400 301 401
rect 302 400 303 401
rect 303 400 304 401
rect 305 400 306 401
rect 300 401 306 405
rect 300 405 301 406
rect 302 405 303 406
rect 303 405 304 406
rect 305 405 306 406
rect 300 160 301 161
rect 302 160 303 161
rect 303 160 304 161
rect 305 160 306 161
rect 300 161 306 165
rect 300 165 301 166
rect 302 165 303 166
rect 303 165 304 166
rect 305 165 306 166
rect 0 220 1 221
rect 2 220 3 221
rect 3 220 4 221
rect 5 220 6 221
rect 0 221 6 225
rect 0 225 1 226
rect 2 225 3 226
rect 3 225 4 226
rect 5 225 6 226
rect 380 140 381 141
rect 382 140 383 141
rect 383 140 384 141
rect 385 140 386 141
rect 380 141 386 145
rect 380 145 381 146
rect 382 145 383 146
rect 383 145 384 146
rect 385 145 386 146
rect 80 40 81 41
rect 82 40 83 41
rect 83 40 84 41
rect 85 40 86 41
rect 80 41 86 45
rect 80 45 81 46
rect 82 45 83 46
rect 83 45 84 46
rect 85 45 86 46
rect 120 340 121 341
rect 122 340 123 341
rect 123 340 124 341
rect 125 340 126 341
rect 120 341 126 345
rect 120 345 121 346
rect 122 345 123 346
rect 123 345 124 346
rect 125 345 126 346
rect 60 300 61 301
rect 62 300 63 301
rect 63 300 64 301
rect 65 300 66 301
rect 60 301 66 305
rect 60 305 61 306
rect 62 305 63 306
rect 63 305 64 306
rect 65 305 66 306
rect 240 0 241 1
rect 242 0 243 1
rect 243 0 244 1
rect 245 0 246 1
rect 240 1 246 5
rect 240 5 241 6
rect 242 5 243 6
rect 243 5 244 6
rect 245 5 246 6
rect 280 240 281 241
rect 282 240 283 241
rect 283 240 284 241
rect 285 240 286 241
rect 280 241 286 245
rect 280 245 281 246
rect 282 245 283 246
rect 283 245 284 246
rect 285 245 286 246
rect 40 320 41 321
rect 42 320 43 321
rect 43 320 44 321
rect 45 320 46 321
rect 40 321 46 325
rect 40 325 41 326
rect 42 325 43 326
rect 43 325 44 326
rect 45 325 46 326
rect 200 100 201 101
rect 202 100 203 101
rect 203 100 204 101
rect 205 100 206 101
rect 200 101 206 105
rect 200 105 201 106
rect 202 105 203 106
rect 203 105 204 106
rect 205 105 206 106
rect 300 100 301 101
rect 302 100 303 101
rect 303 100 304 101
rect 305 100 306 101
rect 300 101 306 105
rect 300 105 301 106
rect 302 105 303 106
rect 303 105 304 106
rect 305 105 306 106
rect 320 300 321 301
rect 322 300 323 301
rect 323 300 324 301
rect 325 300 326 301
rect 320 301 326 305
rect 320 305 321 306
rect 322 305 323 306
rect 323 305 324 306
rect 325 305 326 306
rect 0 120 1 121
rect 2 120 3 121
rect 3 120 4 121
rect 5 120 6 121
rect 0 121 6 125
rect 0 125 1 126
rect 2 125 3 126
rect 3 125 4 126
rect 5 125 6 126
rect 420 240 421 241
rect 422 240 423 241
rect 423 240 424 241
rect 425 240 426 241
rect 420 241 426 245
rect 420 245 421 246
rect 422 245 423 246
rect 423 245 424 246
rect 425 245 426 246
rect 300 340 301 341
rect 302 340 303 341
rect 303 340 304 341
rect 305 340 306 341
rect 300 341 306 345
rect 300 345 301 346
rect 302 345 303 346
rect 303 345 304 346
rect 305 345 306 346
rect 160 200 161 201
rect 162 200 163 201
rect 163 200 164 201
rect 165 200 166 201
rect 160 201 166 205
rect 160 205 161 206
rect 162 205 163 206
rect 163 205 164 206
rect 165 205 166 206
rect 100 140 101 141
rect 102 140 103 141
rect 103 140 104 141
rect 105 140 106 141
rect 100 141 106 145
rect 100 145 101 146
rect 102 145 103 146
rect 103 145 104 146
rect 105 145 106 146
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect 380 280 381 281
rect 382 280 383 281
rect 383 280 384 281
rect 385 280 386 281
rect 380 281 386 285
rect 380 285 381 286
rect 382 285 383 286
rect 383 285 384 286
rect 385 285 386 286
rect 20 160 21 161
rect 22 160 23 161
rect 23 160 24 161
rect 25 160 26 161
rect 20 161 26 165
rect 20 165 21 166
rect 22 165 23 166
rect 23 165 24 166
rect 25 165 26 166
rect 120 180 121 181
rect 122 180 123 181
rect 123 180 124 181
rect 125 180 126 181
rect 120 181 126 185
rect 120 185 121 186
rect 122 185 123 186
rect 123 185 124 186
rect 125 185 126 186
rect 120 120 121 121
rect 122 120 123 121
rect 123 120 124 121
rect 125 120 126 121
rect 120 121 126 125
rect 120 125 121 126
rect 122 125 123 126
rect 123 125 124 126
rect 125 125 126 126
rect 420 200 421 201
rect 422 200 423 201
rect 423 200 424 201
rect 425 200 426 201
rect 420 201 426 205
rect 420 205 421 206
rect 422 205 423 206
rect 423 205 424 206
rect 425 205 426 206
rect 220 240 221 241
rect 222 240 223 241
rect 223 240 224 241
rect 225 240 226 241
rect 220 241 226 245
rect 220 245 221 246
rect 222 245 223 246
rect 223 245 224 246
rect 225 245 226 246
rect 240 240 241 241
rect 242 240 243 241
rect 243 240 244 241
rect 245 240 246 241
rect 240 241 246 245
rect 240 245 241 246
rect 242 245 243 246
rect 243 245 244 246
rect 245 245 246 246
rect 420 220 421 221
rect 422 220 423 221
rect 423 220 424 221
rect 425 220 426 221
rect 420 221 426 225
rect 420 225 421 226
rect 422 225 423 226
rect 423 225 424 226
rect 425 225 426 226
rect 180 420 181 421
rect 182 420 183 421
rect 183 420 184 421
rect 185 420 186 421
rect 180 421 186 425
rect 180 425 181 426
rect 182 425 183 426
rect 183 425 184 426
rect 185 425 186 426
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect 340 400 341 401
rect 342 400 343 401
rect 343 400 344 401
rect 345 400 346 401
rect 340 401 346 405
rect 340 405 341 406
rect 342 405 343 406
rect 343 405 344 406
rect 345 405 346 406
rect 80 220 81 221
rect 82 220 83 221
rect 83 220 84 221
rect 85 220 86 221
rect 80 221 86 225
rect 80 225 81 226
rect 82 225 83 226
rect 83 225 84 226
rect 85 225 86 226
rect 40 240 41 241
rect 42 240 43 241
rect 43 240 44 241
rect 45 240 46 241
rect 40 241 46 245
rect 40 245 41 246
rect 42 245 43 246
rect 43 245 44 246
rect 45 245 46 246
rect 180 360 181 361
rect 182 360 183 361
rect 183 360 184 361
rect 185 360 186 361
rect 180 361 186 365
rect 180 365 181 366
rect 182 365 183 366
rect 183 365 184 366
rect 185 365 186 366
rect 340 220 341 221
rect 342 220 343 221
rect 343 220 344 221
rect 345 220 346 221
rect 340 221 346 225
rect 340 225 341 226
rect 342 225 343 226
rect 343 225 344 226
rect 345 225 346 226
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect 280 0 281 1
rect 282 0 283 1
rect 283 0 284 1
rect 285 0 286 1
rect 280 1 286 5
rect 280 5 281 6
rect 282 5 283 6
rect 283 5 284 6
rect 285 5 286 6
rect 260 160 261 161
rect 262 160 263 161
rect 263 160 264 161
rect 265 160 266 161
rect 260 161 266 165
rect 260 165 261 166
rect 262 165 263 166
rect 263 165 264 166
rect 265 165 266 166
rect 280 320 281 321
rect 282 320 283 321
rect 283 320 284 321
rect 285 320 286 321
rect 280 321 286 325
rect 280 325 281 326
rect 282 325 283 326
rect 283 325 284 326
rect 285 325 286 326
rect 120 220 121 221
rect 122 220 123 221
rect 123 220 124 221
rect 125 220 126 221
rect 120 221 126 225
rect 120 225 121 226
rect 122 225 123 226
rect 123 225 124 226
rect 125 225 126 226
rect 60 160 61 161
rect 62 160 63 161
rect 63 160 64 161
rect 65 160 66 161
rect 60 161 66 165
rect 60 165 61 166
rect 62 165 63 166
rect 63 165 64 166
rect 65 165 66 166
rect 260 120 261 121
rect 262 120 263 121
rect 263 120 264 121
rect 265 120 266 121
rect 260 121 266 125
rect 260 125 261 126
rect 262 125 263 126
rect 263 125 264 126
rect 265 125 266 126
rect 160 100 161 101
rect 162 100 163 101
rect 163 100 164 101
rect 165 100 166 101
rect 160 101 166 105
rect 160 105 161 106
rect 162 105 163 106
rect 163 105 164 106
rect 165 105 166 106
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect 360 220 361 221
rect 362 220 363 221
rect 363 220 364 221
rect 365 220 366 221
rect 360 221 366 225
rect 360 225 361 226
rect 362 225 363 226
rect 363 225 364 226
rect 365 225 366 226
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect 100 400 101 401
rect 102 400 103 401
rect 103 400 104 401
rect 105 400 106 401
rect 100 401 106 405
rect 100 405 101 406
rect 102 405 103 406
rect 103 405 104 406
rect 105 405 106 406
rect 420 120 421 121
rect 422 120 423 121
rect 423 120 424 121
rect 425 120 426 121
rect 420 121 426 125
rect 420 125 421 126
rect 422 125 423 126
rect 423 125 424 126
rect 425 125 426 126
rect 20 180 21 181
rect 22 180 23 181
rect 23 180 24 181
rect 25 180 26 181
rect 20 181 26 185
rect 20 185 21 186
rect 22 185 23 186
rect 23 185 24 186
rect 25 185 26 186
rect 200 60 201 61
rect 202 60 203 61
rect 203 60 204 61
rect 205 60 206 61
rect 200 61 206 65
rect 200 65 201 66
rect 202 65 203 66
rect 203 65 204 66
rect 205 65 206 66
rect 80 80 81 81
rect 82 80 83 81
rect 83 80 84 81
rect 85 80 86 81
rect 80 81 86 85
rect 80 85 81 86
rect 82 85 83 86
rect 83 85 84 86
rect 85 85 86 86
rect 240 400 241 401
rect 242 400 243 401
rect 243 400 244 401
rect 245 400 246 401
rect 240 401 246 405
rect 240 405 241 406
rect 242 405 243 406
rect 243 405 244 406
rect 245 405 246 406
rect 60 240 61 241
rect 62 240 63 241
rect 63 240 64 241
rect 65 240 66 241
rect 60 241 66 245
rect 60 245 61 246
rect 62 245 63 246
rect 63 245 64 246
rect 65 245 66 246
rect 140 160 141 161
rect 142 160 143 161
rect 143 160 144 161
rect 145 160 146 161
rect 140 161 146 165
rect 140 165 141 166
rect 142 165 143 166
rect 143 165 144 166
rect 145 165 146 166
rect 300 320 301 321
rect 302 320 303 321
rect 303 320 304 321
rect 305 320 306 321
rect 300 321 306 325
rect 300 325 301 326
rect 302 325 303 326
rect 303 325 304 326
rect 305 325 306 326
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect 200 20 201 21
rect 202 20 203 21
rect 203 20 204 21
rect 205 20 206 21
rect 200 21 206 25
rect 200 25 201 26
rect 202 25 203 26
rect 203 25 204 26
rect 205 25 206 26
rect 280 20 281 21
rect 282 20 283 21
rect 283 20 284 21
rect 285 20 286 21
rect 280 21 286 25
rect 280 25 281 26
rect 282 25 283 26
rect 283 25 284 26
rect 285 25 286 26
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect 180 320 181 321
rect 182 320 183 321
rect 183 320 184 321
rect 185 320 186 321
rect 180 321 186 325
rect 180 325 181 326
rect 182 325 183 326
rect 183 325 184 326
rect 185 325 186 326
rect 220 140 221 141
rect 222 140 223 141
rect 223 140 224 141
rect 225 140 226 141
rect 220 141 226 145
rect 220 145 221 146
rect 222 145 223 146
rect 223 145 224 146
rect 225 145 226 146
rect 320 60 321 61
rect 322 60 323 61
rect 323 60 324 61
rect 325 60 326 61
rect 320 61 326 65
rect 320 65 321 66
rect 322 65 323 66
rect 323 65 324 66
rect 325 65 326 66
rect 20 220 21 221
rect 22 220 23 221
rect 23 220 24 221
rect 25 220 26 221
rect 20 221 26 225
rect 20 225 21 226
rect 22 225 23 226
rect 23 225 24 226
rect 25 225 26 226
rect 280 260 281 261
rect 282 260 283 261
rect 283 260 284 261
rect 285 260 286 261
rect 280 261 286 265
rect 280 265 281 266
rect 282 265 283 266
rect 283 265 284 266
rect 285 265 286 266
rect 140 280 141 281
rect 142 280 143 281
rect 143 280 144 281
rect 145 280 146 281
rect 140 281 146 285
rect 140 285 141 286
rect 142 285 143 286
rect 143 285 144 286
rect 145 285 146 286
rect 300 280 301 281
rect 302 280 303 281
rect 303 280 304 281
rect 305 280 306 281
rect 300 281 306 285
rect 300 285 301 286
rect 302 285 303 286
rect 303 285 304 286
rect 305 285 306 286
rect 400 180 401 181
rect 402 180 403 181
rect 403 180 404 181
rect 405 180 406 181
rect 400 181 406 185
rect 400 185 401 186
rect 402 185 403 186
rect 403 185 404 186
rect 405 185 406 186
rect 140 120 141 121
rect 142 120 143 121
rect 143 120 144 121
rect 145 120 146 121
rect 140 121 146 125
rect 140 125 141 126
rect 142 125 143 126
rect 143 125 144 126
rect 145 125 146 126
rect 120 140 121 141
rect 122 140 123 141
rect 123 140 124 141
rect 125 140 126 141
rect 120 141 126 145
rect 120 145 121 146
rect 122 145 123 146
rect 123 145 124 146
rect 125 145 126 146
rect 260 200 261 201
rect 262 200 263 201
rect 263 200 264 201
rect 265 200 266 201
rect 260 201 266 205
rect 260 205 261 206
rect 262 205 263 206
rect 263 205 264 206
rect 265 205 266 206
rect 160 220 161 221
rect 162 220 163 221
rect 163 220 164 221
rect 165 220 166 221
rect 160 221 166 225
rect 160 225 161 226
rect 162 225 163 226
rect 163 225 164 226
rect 165 225 166 226
rect 260 460 261 461
rect 262 460 263 461
rect 263 460 264 461
rect 265 460 266 461
rect 260 461 266 465
rect 260 465 261 466
rect 262 465 263 466
rect 263 465 264 466
rect 265 465 266 466
rect 120 60 121 61
rect 122 60 123 61
rect 123 60 124 61
rect 125 60 126 61
rect 120 61 126 65
rect 120 65 121 66
rect 122 65 123 66
rect 123 65 124 66
rect 125 65 126 66
rect 300 360 301 361
rect 302 360 303 361
rect 303 360 304 361
rect 305 360 306 361
rect 300 361 306 365
rect 300 365 301 366
rect 302 365 303 366
rect 303 365 304 366
rect 305 365 306 366
rect 200 140 201 141
rect 202 140 203 141
rect 203 140 204 141
rect 205 140 206 141
rect 200 141 206 145
rect 200 145 201 146
rect 202 145 203 146
rect 203 145 204 146
rect 205 145 206 146
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect 100 160 101 161
rect 102 160 103 161
rect 103 160 104 161
rect 105 160 106 161
rect 100 161 106 165
rect 100 165 101 166
rect 102 165 103 166
rect 103 165 104 166
rect 105 165 106 166
rect 240 40 241 41
rect 242 40 243 41
rect 243 40 244 41
rect 245 40 246 41
rect 240 41 246 45
rect 240 45 241 46
rect 242 45 243 46
rect 243 45 244 46
rect 245 45 246 46
rect 220 300 221 301
rect 222 300 223 301
rect 223 300 224 301
rect 225 300 226 301
rect 220 301 226 305
rect 220 305 221 306
rect 222 305 223 306
rect 223 305 224 306
rect 225 305 226 306
rect 200 80 201 81
rect 202 80 203 81
rect 203 80 204 81
rect 205 80 206 81
rect 200 81 206 85
rect 200 85 201 86
rect 202 85 203 86
rect 203 85 204 86
rect 205 85 206 86
rect 200 40 201 41
rect 202 40 203 41
rect 203 40 204 41
rect 205 40 206 41
rect 200 41 206 45
rect 200 45 201 46
rect 202 45 203 46
rect 203 45 204 46
rect 205 45 206 46
rect 320 360 321 361
rect 322 360 323 361
rect 323 360 324 361
rect 325 360 326 361
rect 320 361 326 365
rect 320 365 321 366
rect 322 365 323 366
rect 323 365 324 366
rect 325 365 326 366
rect 340 280 341 281
rect 342 280 343 281
rect 343 280 344 281
rect 345 280 346 281
rect 340 281 346 285
rect 340 285 341 286
rect 342 285 343 286
rect 343 285 344 286
rect 345 285 346 286
rect 360 100 361 101
rect 362 100 363 101
rect 363 100 364 101
rect 365 100 366 101
rect 360 101 366 105
rect 360 105 361 106
rect 362 105 363 106
rect 363 105 364 106
rect 365 105 366 106
rect 80 140 81 141
rect 82 140 83 141
rect 83 140 84 141
rect 85 140 86 141
rect 80 141 86 145
rect 80 145 81 146
rect 82 145 83 146
rect 83 145 84 146
rect 85 145 86 146
rect 60 80 61 81
rect 62 80 63 81
rect 63 80 64 81
rect 65 80 66 81
rect 60 81 66 85
rect 60 85 61 86
rect 62 85 63 86
rect 63 85 64 86
rect 65 85 66 86
rect 120 280 121 281
rect 122 280 123 281
rect 123 280 124 281
rect 125 280 126 281
rect 120 281 126 285
rect 120 285 121 286
rect 122 285 123 286
rect 123 285 124 286
rect 125 285 126 286
rect 260 240 261 241
rect 262 240 263 241
rect 263 240 264 241
rect 265 240 266 241
rect 260 241 266 245
rect 260 245 261 246
rect 262 245 263 246
rect 263 245 264 246
rect 265 245 266 246
rect 320 380 321 381
rect 322 380 323 381
rect 323 380 324 381
rect 325 380 326 381
rect 320 381 326 385
rect 320 385 321 386
rect 322 385 323 386
rect 323 385 324 386
rect 325 385 326 386
rect 160 360 161 361
rect 162 360 163 361
rect 163 360 164 361
rect 165 360 166 361
rect 160 361 166 365
rect 160 365 161 366
rect 162 365 163 366
rect 163 365 164 366
rect 165 365 166 366
rect 220 100 221 101
rect 222 100 223 101
rect 223 100 224 101
rect 225 100 226 101
rect 220 101 226 105
rect 220 105 221 106
rect 222 105 223 106
rect 223 105 224 106
rect 225 105 226 106
rect 180 80 181 81
rect 182 80 183 81
rect 183 80 184 81
rect 185 80 186 81
rect 180 81 186 85
rect 180 85 181 86
rect 182 85 183 86
rect 183 85 184 86
rect 185 85 186 86
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect 240 320 241 321
rect 242 320 243 321
rect 243 320 244 321
rect 245 320 246 321
rect 240 321 246 325
rect 240 325 241 326
rect 242 325 243 326
rect 243 325 244 326
rect 245 325 246 326
rect 300 300 301 301
rect 302 300 303 301
rect 303 300 304 301
rect 305 300 306 301
rect 300 301 306 305
rect 300 305 301 306
rect 302 305 303 306
rect 303 305 304 306
rect 305 305 306 306
rect 200 320 201 321
rect 202 320 203 321
rect 203 320 204 321
rect 205 320 206 321
rect 200 321 206 325
rect 200 325 201 326
rect 202 325 203 326
rect 203 325 204 326
rect 205 325 206 326
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect 60 320 61 321
rect 62 320 63 321
rect 63 320 64 321
rect 65 320 66 321
rect 60 321 66 325
rect 60 325 61 326
rect 62 325 63 326
rect 63 325 64 326
rect 65 325 66 326
rect 220 160 221 161
rect 222 160 223 161
rect 223 160 224 161
rect 225 160 226 161
rect 220 161 226 165
rect 220 165 221 166
rect 222 165 223 166
rect 223 165 224 166
rect 225 165 226 166
rect 80 380 81 381
rect 82 380 83 381
rect 83 380 84 381
rect 85 380 86 381
rect 80 381 86 385
rect 80 385 81 386
rect 82 385 83 386
rect 83 385 84 386
rect 85 385 86 386
rect 260 380 261 381
rect 262 380 263 381
rect 263 380 264 381
rect 265 380 266 381
rect 260 381 266 385
rect 260 385 261 386
rect 262 385 263 386
rect 263 385 264 386
rect 265 385 266 386
rect 340 340 341 341
rect 342 340 343 341
rect 343 340 344 341
rect 345 340 346 341
rect 340 341 346 345
rect 340 345 341 346
rect 342 345 343 346
rect 343 345 344 346
rect 345 345 346 346
rect 280 160 281 161
rect 282 160 283 161
rect 283 160 284 161
rect 285 160 286 161
rect 280 161 286 165
rect 280 165 281 166
rect 282 165 283 166
rect 283 165 284 166
rect 285 165 286 166
rect 20 280 21 281
rect 22 280 23 281
rect 23 280 24 281
rect 25 280 26 281
rect 20 281 26 285
rect 20 285 21 286
rect 22 285 23 286
rect 23 285 24 286
rect 25 285 26 286
rect 360 280 361 281
rect 362 280 363 281
rect 363 280 364 281
rect 365 280 366 281
rect 360 281 366 285
rect 360 285 361 286
rect 362 285 363 286
rect 363 285 364 286
rect 365 285 366 286
rect 40 220 41 221
rect 42 220 43 221
rect 43 220 44 221
rect 45 220 46 221
rect 40 221 46 225
rect 40 225 41 226
rect 42 225 43 226
rect 43 225 44 226
rect 45 225 46 226
rect 140 60 141 61
rect 142 60 143 61
rect 143 60 144 61
rect 145 60 146 61
rect 140 61 146 65
rect 140 65 141 66
rect 142 65 143 66
rect 143 65 144 66
rect 145 65 146 66
rect 180 160 181 161
rect 182 160 183 161
rect 183 160 184 161
rect 185 160 186 161
rect 180 161 186 165
rect 180 165 181 166
rect 182 165 183 166
rect 183 165 184 166
rect 185 165 186 166
rect 360 380 361 381
rect 362 380 363 381
rect 363 380 364 381
rect 365 380 366 381
rect 360 381 366 385
rect 360 385 361 386
rect 362 385 363 386
rect 363 385 364 386
rect 365 385 366 386
rect 80 180 81 181
rect 82 180 83 181
rect 83 180 84 181
rect 85 180 86 181
rect 80 181 86 185
rect 80 185 81 186
rect 82 185 83 186
rect 83 185 84 186
rect 85 185 86 186
rect 220 260 221 261
rect 222 260 223 261
rect 223 260 224 261
rect 225 260 226 261
rect 220 261 226 265
rect 220 265 221 266
rect 222 265 223 266
rect 223 265 224 266
rect 225 265 226 266
rect 340 140 341 141
rect 342 140 343 141
rect 343 140 344 141
rect 345 140 346 141
rect 340 141 346 145
rect 340 145 341 146
rect 342 145 343 146
rect 343 145 344 146
rect 345 145 346 146
rect 140 40 141 41
rect 142 40 143 41
rect 143 40 144 41
rect 145 40 146 41
rect 140 41 146 45
rect 140 45 141 46
rect 142 45 143 46
rect 143 45 144 46
rect 145 45 146 46
rect 100 380 101 381
rect 102 380 103 381
rect 103 380 104 381
rect 105 380 106 381
rect 100 381 106 385
rect 100 385 101 386
rect 102 385 103 386
rect 103 385 104 386
rect 105 385 106 386
rect 340 200 341 201
rect 342 200 343 201
rect 343 200 344 201
rect 345 200 346 201
rect 340 201 346 205
rect 340 205 341 206
rect 342 205 343 206
rect 343 205 344 206
rect 345 205 346 206
rect 320 280 321 281
rect 322 280 323 281
rect 323 280 324 281
rect 325 280 326 281
rect 320 281 326 285
rect 320 285 321 286
rect 322 285 323 286
rect 323 285 324 286
rect 325 285 326 286
rect 200 260 201 261
rect 202 260 203 261
rect 203 260 204 261
rect 205 260 206 261
rect 200 261 206 265
rect 200 265 201 266
rect 202 265 203 266
rect 203 265 204 266
rect 205 265 206 266
rect 200 400 201 401
rect 202 400 203 401
rect 203 400 204 401
rect 205 400 206 401
rect 200 401 206 405
rect 200 405 201 406
rect 202 405 203 406
rect 203 405 204 406
rect 205 405 206 406
rect 80 100 81 101
rect 82 100 83 101
rect 83 100 84 101
rect 85 100 86 101
rect 80 101 86 105
rect 80 105 81 106
rect 82 105 83 106
rect 83 105 84 106
rect 85 105 86 106
rect 60 100 61 101
rect 62 100 63 101
rect 63 100 64 101
rect 65 100 66 101
rect 60 101 66 105
rect 60 105 61 106
rect 62 105 63 106
rect 63 105 64 106
rect 65 105 66 106
rect 140 80 141 81
rect 142 80 143 81
rect 143 80 144 81
rect 145 80 146 81
rect 140 81 146 85
rect 140 85 141 86
rect 142 85 143 86
rect 143 85 144 86
rect 145 85 146 86
rect 280 140 281 141
rect 282 140 283 141
rect 283 140 284 141
rect 285 140 286 141
rect 280 141 286 145
rect 280 145 281 146
rect 282 145 283 146
rect 283 145 284 146
rect 285 145 286 146
rect 300 180 301 181
rect 302 180 303 181
rect 303 180 304 181
rect 305 180 306 181
rect 300 181 306 185
rect 300 185 301 186
rect 302 185 303 186
rect 303 185 304 186
rect 305 185 306 186
rect 340 300 341 301
rect 342 300 343 301
rect 343 300 344 301
rect 345 300 346 301
rect 340 301 346 305
rect 340 305 341 306
rect 342 305 343 306
rect 343 305 344 306
rect 345 305 346 306
rect 400 300 401 301
rect 402 300 403 301
rect 403 300 404 301
rect 405 300 406 301
rect 400 301 406 305
rect 400 305 401 306
rect 402 305 403 306
rect 403 305 404 306
rect 405 305 406 306
rect 220 360 221 361
rect 222 360 223 361
rect 223 360 224 361
rect 225 360 226 361
rect 220 361 226 365
rect 220 365 221 366
rect 222 365 223 366
rect 223 365 224 366
rect 225 365 226 366
rect 180 220 181 221
rect 182 220 183 221
rect 183 220 184 221
rect 185 220 186 221
rect 180 221 186 225
rect 180 225 181 226
rect 182 225 183 226
rect 183 225 184 226
rect 185 225 186 226
rect 160 60 161 61
rect 162 60 163 61
rect 163 60 164 61
rect 165 60 166 61
rect 160 61 166 65
rect 160 65 161 66
rect 162 65 163 66
rect 163 65 164 66
rect 165 65 166 66
rect 40 180 41 181
rect 42 180 43 181
rect 43 180 44 181
rect 45 180 46 181
rect 40 181 46 185
rect 40 185 41 186
rect 42 185 43 186
rect 43 185 44 186
rect 45 185 46 186
rect 60 280 61 281
rect 62 280 63 281
rect 63 280 64 281
rect 65 280 66 281
rect 60 281 66 285
rect 60 285 61 286
rect 62 285 63 286
rect 63 285 64 286
rect 65 285 66 286
rect 180 180 181 181
rect 182 180 183 181
rect 183 180 184 181
rect 185 180 186 181
rect 180 181 186 185
rect 180 185 181 186
rect 182 185 183 186
rect 183 185 184 186
rect 185 185 186 186
rect 160 120 161 121
rect 162 120 163 121
rect 163 120 164 121
rect 165 120 166 121
rect 160 121 166 125
rect 160 125 161 126
rect 162 125 163 126
rect 163 125 164 126
rect 165 125 166 126
rect 380 320 381 321
rect 382 320 383 321
rect 383 320 384 321
rect 385 320 386 321
rect 380 321 386 325
rect 380 325 381 326
rect 382 325 383 326
rect 383 325 384 326
rect 385 325 386 326
rect 240 200 241 201
rect 242 200 243 201
rect 243 200 244 201
rect 245 200 246 201
rect 240 201 246 205
rect 240 205 241 206
rect 242 205 243 206
rect 243 205 244 206
rect 245 205 246 206
rect 80 340 81 341
rect 82 340 83 341
rect 83 340 84 341
rect 85 340 86 341
rect 80 341 86 345
rect 80 345 81 346
rect 82 345 83 346
rect 83 345 84 346
rect 85 345 86 346
rect 360 300 361 301
rect 362 300 363 301
rect 363 300 364 301
rect 365 300 366 301
rect 360 301 366 305
rect 360 305 361 306
rect 362 305 363 306
rect 363 305 364 306
rect 365 305 366 306
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect 300 380 301 381
rect 302 380 303 381
rect 303 380 304 381
rect 305 380 306 381
rect 300 381 306 385
rect 300 385 301 386
rect 302 385 303 386
rect 303 385 304 386
rect 305 385 306 386
rect 320 260 321 261
rect 322 260 323 261
rect 323 260 324 261
rect 325 260 326 261
rect 320 261 326 265
rect 320 265 321 266
rect 322 265 323 266
rect 323 265 324 266
rect 325 265 326 266
rect 340 240 341 241
rect 342 240 343 241
rect 343 240 344 241
rect 345 240 346 241
rect 340 241 346 245
rect 340 245 341 246
rect 342 245 343 246
rect 343 245 344 246
rect 345 245 346 246
rect 120 160 121 161
rect 122 160 123 161
rect 123 160 124 161
rect 125 160 126 161
rect 120 161 126 165
rect 120 165 121 166
rect 122 165 123 166
rect 123 165 124 166
rect 125 165 126 166
rect 280 180 281 181
rect 282 180 283 181
rect 283 180 284 181
rect 285 180 286 181
rect 280 181 286 185
rect 280 185 281 186
rect 282 185 283 186
rect 283 185 284 186
rect 285 185 286 186
rect 220 340 221 341
rect 222 340 223 341
rect 223 340 224 341
rect 225 340 226 341
rect 220 341 226 345
rect 220 345 221 346
rect 222 345 223 346
rect 223 345 224 346
rect 225 345 226 346
rect 100 220 101 221
rect 102 220 103 221
rect 103 220 104 221
rect 105 220 106 221
rect 100 221 106 225
rect 100 225 101 226
rect 102 225 103 226
rect 103 225 104 226
rect 105 225 106 226
rect 180 140 181 141
rect 182 140 183 141
rect 183 140 184 141
rect 185 140 186 141
rect 180 141 186 145
rect 180 145 181 146
rect 182 145 183 146
rect 183 145 184 146
rect 185 145 186 146
rect 360 340 361 341
rect 362 340 363 341
rect 363 340 364 341
rect 365 340 366 341
rect 360 341 366 345
rect 360 345 361 346
rect 362 345 363 346
rect 363 345 364 346
rect 365 345 366 346
rect 60 220 61 221
rect 62 220 63 221
rect 63 220 64 221
rect 65 220 66 221
rect 60 221 66 225
rect 60 225 61 226
rect 62 225 63 226
rect 63 225 64 226
rect 65 225 66 226
rect 280 280 281 281
rect 282 280 283 281
rect 283 280 284 281
rect 285 280 286 281
rect 280 281 286 285
rect 280 285 281 286
rect 282 285 283 286
rect 283 285 284 286
rect 285 285 286 286
rect 320 100 321 101
rect 322 100 323 101
rect 323 100 324 101
rect 325 100 326 101
rect 320 101 326 105
rect 320 105 321 106
rect 322 105 323 106
rect 323 105 324 106
rect 325 105 326 106
rect 380 220 381 221
rect 382 220 383 221
rect 383 220 384 221
rect 385 220 386 221
rect 380 221 386 225
rect 380 225 381 226
rect 382 225 383 226
rect 383 225 384 226
rect 385 225 386 226
rect 120 80 121 81
rect 122 80 123 81
rect 123 80 124 81
rect 125 80 126 81
rect 120 81 126 85
rect 120 85 121 86
rect 122 85 123 86
rect 123 85 124 86
rect 125 85 126 86
rect 320 140 321 141
rect 322 140 323 141
rect 323 140 324 141
rect 325 140 326 141
rect 320 141 326 145
rect 320 145 321 146
rect 322 145 323 146
rect 323 145 324 146
rect 325 145 326 146
rect 0 260 1 261
rect 2 260 3 261
rect 3 260 4 261
rect 5 260 6 261
rect 0 261 6 265
rect 0 265 1 266
rect 2 265 3 266
rect 3 265 4 266
rect 5 265 6 266
rect 320 40 321 41
rect 322 40 323 41
rect 323 40 324 41
rect 325 40 326 41
rect 320 41 326 45
rect 320 45 321 46
rect 322 45 323 46
rect 323 45 324 46
rect 325 45 326 46
rect 220 220 221 221
rect 222 220 223 221
rect 223 220 224 221
rect 225 220 226 221
rect 220 221 226 225
rect 220 225 221 226
rect 222 225 223 226
rect 223 225 224 226
rect 225 225 226 226
rect 100 300 101 301
rect 102 300 103 301
rect 103 300 104 301
rect 105 300 106 301
rect 100 301 106 305
rect 100 305 101 306
rect 102 305 103 306
rect 103 305 104 306
rect 105 305 106 306
rect 280 80 281 81
rect 282 80 283 81
rect 283 80 284 81
rect 285 80 286 81
rect 280 81 286 85
rect 280 85 281 86
rect 282 85 283 86
rect 283 85 284 86
rect 285 85 286 86
rect 180 20 181 21
rect 182 20 183 21
rect 183 20 184 21
rect 185 20 186 21
rect 180 21 186 25
rect 180 25 181 26
rect 182 25 183 26
rect 183 25 184 26
rect 185 25 186 26
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect 220 60 221 61
rect 222 60 223 61
rect 223 60 224 61
rect 225 60 226 61
rect 220 61 226 65
rect 220 65 221 66
rect 222 65 223 66
rect 223 65 224 66
rect 225 65 226 66
rect 200 200 201 201
rect 202 200 203 201
rect 203 200 204 201
rect 205 200 206 201
rect 200 201 206 205
rect 200 205 201 206
rect 202 205 203 206
rect 203 205 204 206
rect 205 205 206 206
rect 260 140 261 141
rect 262 140 263 141
rect 263 140 264 141
rect 265 140 266 141
rect 260 141 266 145
rect 260 145 261 146
rect 262 145 263 146
rect 263 145 264 146
rect 265 145 266 146
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect 280 200 281 201
rect 282 200 283 201
rect 283 200 284 201
rect 285 200 286 201
rect 280 201 286 205
rect 280 205 281 206
rect 282 205 283 206
rect 283 205 284 206
rect 285 205 286 206
rect 300 220 301 221
rect 302 220 303 221
rect 303 220 304 221
rect 305 220 306 221
rect 300 221 306 225
rect 300 225 301 226
rect 302 225 303 226
rect 303 225 304 226
rect 305 225 306 226
rect 220 180 221 181
rect 222 180 223 181
rect 223 180 224 181
rect 225 180 226 181
rect 220 181 226 185
rect 220 185 221 186
rect 222 185 223 186
rect 223 185 224 186
rect 225 185 226 186
rect 240 360 241 361
rect 242 360 243 361
rect 243 360 244 361
rect 245 360 246 361
rect 240 361 246 365
rect 240 365 241 366
rect 242 365 243 366
rect 243 365 244 366
rect 245 365 246 366
rect 440 200 441 201
rect 442 200 443 201
rect 443 200 444 201
rect 445 200 446 201
rect 440 201 446 205
rect 440 205 441 206
rect 442 205 443 206
rect 443 205 444 206
rect 445 205 446 206
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect 160 20 161 21
rect 162 20 163 21
rect 163 20 164 21
rect 165 20 166 21
rect 160 21 166 25
rect 160 25 161 26
rect 162 25 163 26
rect 163 25 164 26
rect 165 25 166 26
rect 160 80 161 81
rect 162 80 163 81
rect 163 80 164 81
rect 165 80 166 81
rect 160 81 166 85
rect 160 85 161 86
rect 162 85 163 86
rect 163 85 164 86
rect 165 85 166 86
rect 160 280 161 281
rect 162 280 163 281
rect 163 280 164 281
rect 165 280 166 281
rect 160 281 166 285
rect 160 285 161 286
rect 162 285 163 286
rect 163 285 164 286
rect 165 285 166 286
rect 40 200 41 201
rect 42 200 43 201
rect 43 200 44 201
rect 45 200 46 201
rect 40 201 46 205
rect 40 205 41 206
rect 42 205 43 206
rect 43 205 44 206
rect 45 205 46 206
rect 200 180 201 181
rect 202 180 203 181
rect 203 180 204 181
rect 205 180 206 181
rect 200 181 206 185
rect 200 185 201 186
rect 202 185 203 186
rect 203 185 204 186
rect 205 185 206 186
rect 180 340 181 341
rect 182 340 183 341
rect 183 340 184 341
rect 185 340 186 341
rect 180 341 186 345
rect 180 345 181 346
rect 182 345 183 346
rect 183 345 184 346
rect 185 345 186 346
rect 80 200 81 201
rect 82 200 83 201
rect 83 200 84 201
rect 85 200 86 201
rect 80 201 86 205
rect 80 205 81 206
rect 82 205 83 206
rect 83 205 84 206
rect 85 205 86 206
rect 300 260 301 261
rect 302 260 303 261
rect 303 260 304 261
rect 305 260 306 261
rect 300 261 306 265
rect 300 265 301 266
rect 302 265 303 266
rect 303 265 304 266
rect 305 265 306 266
rect 200 380 201 381
rect 202 380 203 381
rect 203 380 204 381
rect 205 380 206 381
rect 200 381 206 385
rect 200 385 201 386
rect 202 385 203 386
rect 203 385 204 386
rect 205 385 206 386
rect 220 280 221 281
rect 222 280 223 281
rect 223 280 224 281
rect 225 280 226 281
rect 220 281 226 285
rect 220 285 221 286
rect 222 285 223 286
rect 223 285 224 286
rect 225 285 226 286
rect 260 420 261 421
rect 262 420 263 421
rect 263 420 264 421
rect 265 420 266 421
rect 260 421 266 425
rect 260 425 261 426
rect 262 425 263 426
rect 263 425 264 426
rect 265 425 266 426
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect 60 340 61 341
rect 62 340 63 341
rect 63 340 64 341
rect 65 340 66 341
rect 60 341 66 345
rect 60 345 61 346
rect 62 345 63 346
rect 63 345 64 346
rect 65 345 66 346
rect 120 260 121 261
rect 122 260 123 261
rect 123 260 124 261
rect 125 260 126 261
rect 120 261 126 265
rect 120 265 121 266
rect 122 265 123 266
rect 123 265 124 266
rect 125 265 126 266
rect 140 100 141 101
rect 142 100 143 101
rect 143 100 144 101
rect 145 100 146 101
rect 140 101 146 105
rect 140 105 141 106
rect 142 105 143 106
rect 143 105 144 106
rect 145 105 146 106
rect 340 320 341 321
rect 342 320 343 321
rect 343 320 344 321
rect 345 320 346 321
rect 340 321 346 325
rect 340 325 341 326
rect 342 325 343 326
rect 343 325 344 326
rect 345 325 346 326
rect 140 20 141 21
rect 142 20 143 21
rect 143 20 144 21
rect 145 20 146 21
rect 140 21 146 25
rect 140 25 141 26
rect 142 25 143 26
rect 143 25 144 26
rect 145 25 146 26
rect 60 260 61 261
rect 62 260 63 261
rect 63 260 64 261
rect 65 260 66 261
rect 60 261 66 265
rect 60 265 61 266
rect 62 265 63 266
rect 63 265 64 266
rect 65 265 66 266
rect 240 440 241 441
rect 242 440 243 441
rect 243 440 244 441
rect 245 440 246 441
rect 240 441 246 445
rect 240 445 241 446
rect 242 445 243 446
rect 243 445 244 446
rect 245 445 246 446
rect 240 120 241 121
rect 242 120 243 121
rect 243 120 244 121
rect 245 120 246 121
rect 240 121 246 125
rect 240 125 241 126
rect 242 125 243 126
rect 243 125 244 126
rect 245 125 246 126
rect 140 180 141 181
rect 142 180 143 181
rect 143 180 144 181
rect 145 180 146 181
rect 140 181 146 185
rect 140 185 141 186
rect 142 185 143 186
rect 143 185 144 186
rect 145 185 146 186
rect 280 40 281 41
rect 282 40 283 41
rect 283 40 284 41
rect 285 40 286 41
rect 280 41 286 45
rect 280 45 281 46
rect 282 45 283 46
rect 283 45 284 46
rect 285 45 286 46
rect 360 200 361 201
rect 362 200 363 201
rect 363 200 364 201
rect 365 200 366 201
rect 360 201 366 205
rect 360 205 361 206
rect 362 205 363 206
rect 363 205 364 206
rect 365 205 366 206
rect 340 380 341 381
rect 342 380 343 381
rect 343 380 344 381
rect 345 380 346 381
rect 340 381 346 385
rect 340 385 341 386
rect 342 385 343 386
rect 343 385 344 386
rect 345 385 346 386
rect 0 280 1 281
rect 2 280 3 281
rect 3 280 4 281
rect 5 280 6 281
rect 0 281 6 285
rect 0 285 1 286
rect 2 285 3 286
rect 3 285 4 286
rect 5 285 6 286
rect 300 80 301 81
rect 302 80 303 81
rect 303 80 304 81
rect 305 80 306 81
rect 300 81 306 85
rect 300 85 301 86
rect 302 85 303 86
rect 303 85 304 86
rect 305 85 306 86
rect 280 360 281 361
rect 282 360 283 361
rect 283 360 284 361
rect 285 360 286 361
rect 280 361 286 365
rect 280 365 281 366
rect 282 365 283 366
rect 283 365 284 366
rect 285 365 286 366
rect 120 300 121 301
rect 122 300 123 301
rect 123 300 124 301
rect 125 300 126 301
rect 120 301 126 305
rect 120 305 121 306
rect 122 305 123 306
rect 123 305 124 306
rect 125 305 126 306
rect 220 120 221 121
rect 222 120 223 121
rect 223 120 224 121
rect 225 120 226 121
rect 220 121 226 125
rect 220 125 221 126
rect 222 125 223 126
rect 223 125 224 126
rect 225 125 226 126
rect 160 40 161 41
rect 162 40 163 41
rect 163 40 164 41
rect 165 40 166 41
rect 160 41 166 45
rect 160 45 161 46
rect 162 45 163 46
rect 163 45 164 46
rect 165 45 166 46
rect 260 0 261 1
rect 262 0 263 1
rect 263 0 264 1
rect 265 0 266 1
rect 260 1 266 5
rect 260 5 261 6
rect 262 5 263 6
rect 263 5 264 6
rect 265 5 266 6
rect 240 180 241 181
rect 242 180 243 181
rect 243 180 244 181
rect 245 180 246 181
rect 240 181 246 185
rect 240 185 241 186
rect 242 185 243 186
rect 243 185 244 186
rect 245 185 246 186
rect 200 340 201 341
rect 202 340 203 341
rect 203 340 204 341
rect 205 340 206 341
rect 200 341 206 345
rect 200 345 201 346
rect 202 345 203 346
rect 203 345 204 346
rect 205 345 206 346
rect 340 160 341 161
rect 342 160 343 161
rect 343 160 344 161
rect 345 160 346 161
rect 340 161 346 165
rect 340 165 341 166
rect 342 165 343 166
rect 343 165 344 166
rect 345 165 346 166
rect 120 40 121 41
rect 122 40 123 41
rect 123 40 124 41
rect 125 40 126 41
rect 120 41 126 45
rect 120 45 121 46
rect 122 45 123 46
rect 123 45 124 46
rect 125 45 126 46
rect 300 240 301 241
rect 302 240 303 241
rect 303 240 304 241
rect 305 240 306 241
rect 300 241 306 245
rect 300 245 301 246
rect 302 245 303 246
rect 303 245 304 246
rect 305 245 306 246
rect 280 420 281 421
rect 282 420 283 421
rect 283 420 284 421
rect 285 420 286 421
rect 280 421 286 425
rect 280 425 281 426
rect 282 425 283 426
rect 283 425 284 426
rect 285 425 286 426
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect 180 240 181 241
rect 182 240 183 241
rect 183 240 184 241
rect 185 240 186 241
rect 180 241 186 245
rect 180 245 181 246
rect 182 245 183 246
rect 183 245 184 246
rect 185 245 186 246
rect 260 60 261 61
rect 262 60 263 61
rect 263 60 264 61
rect 265 60 266 61
rect 260 61 266 65
rect 260 65 261 66
rect 262 65 263 66
rect 263 65 264 66
rect 265 65 266 66
rect 260 280 261 281
rect 262 280 263 281
rect 263 280 264 281
rect 265 280 266 281
rect 260 281 266 285
rect 260 285 261 286
rect 262 285 263 286
rect 263 285 264 286
rect 265 285 266 286
rect 320 120 321 121
rect 322 120 323 121
rect 323 120 324 121
rect 325 120 326 121
rect 320 121 326 125
rect 320 125 321 126
rect 322 125 323 126
rect 323 125 324 126
rect 325 125 326 126
rect 300 200 301 201
rect 302 200 303 201
rect 303 200 304 201
rect 305 200 306 201
rect 300 201 306 205
rect 300 205 301 206
rect 302 205 303 206
rect 303 205 304 206
rect 305 205 306 206
rect 320 340 321 341
rect 322 340 323 341
rect 323 340 324 341
rect 325 340 326 341
rect 320 341 326 345
rect 320 345 321 346
rect 322 345 323 346
rect 323 345 324 346
rect 325 345 326 346
rect 240 140 241 141
rect 242 140 243 141
rect 243 140 244 141
rect 245 140 246 141
rect 240 141 246 145
rect 240 145 241 146
rect 242 145 243 146
rect 243 145 244 146
rect 245 145 246 146
rect 60 140 61 141
rect 62 140 63 141
rect 63 140 64 141
rect 65 140 66 141
rect 60 141 66 145
rect 60 145 61 146
rect 62 145 63 146
rect 63 145 64 146
rect 65 145 66 146
rect 360 120 361 121
rect 362 120 363 121
rect 363 120 364 121
rect 365 120 366 121
rect 360 121 366 125
rect 360 125 361 126
rect 362 125 363 126
rect 363 125 364 126
rect 365 125 366 126
rect 200 240 201 241
rect 202 240 203 241
rect 203 240 204 241
rect 205 240 206 241
rect 200 241 206 245
rect 200 245 201 246
rect 202 245 203 246
rect 203 245 204 246
rect 205 245 206 246
rect 340 180 341 181
rect 342 180 343 181
rect 343 180 344 181
rect 345 180 346 181
rect 340 181 346 185
rect 340 185 341 186
rect 342 185 343 186
rect 343 185 344 186
rect 345 185 346 186
rect 60 180 61 181
rect 62 180 63 181
rect 63 180 64 181
rect 65 180 66 181
rect 60 181 66 185
rect 60 185 61 186
rect 62 185 63 186
rect 63 185 64 186
rect 65 185 66 186
rect 180 40 181 41
rect 182 40 183 41
rect 183 40 184 41
rect 185 40 186 41
rect 180 41 186 45
rect 180 45 181 46
rect 182 45 183 46
rect 183 45 184 46
rect 185 45 186 46
rect 200 460 201 461
rect 202 460 203 461
rect 203 460 204 461
rect 205 460 206 461
rect 200 461 206 465
rect 200 465 201 466
rect 202 465 203 466
rect 203 465 204 466
rect 205 465 206 466
rect 340 100 341 101
rect 342 100 343 101
rect 343 100 344 101
rect 345 100 346 101
rect 340 101 346 105
rect 340 105 341 106
rect 342 105 343 106
rect 343 105 344 106
rect 345 105 346 106
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect 260 80 261 81
rect 262 80 263 81
rect 263 80 264 81
rect 265 80 266 81
rect 260 81 266 85
rect 260 85 261 86
rect 262 85 263 86
rect 263 85 264 86
rect 265 85 266 86
rect 180 60 181 61
rect 182 60 183 61
rect 183 60 184 61
rect 185 60 186 61
rect 180 61 186 65
rect 180 65 181 66
rect 182 65 183 66
rect 183 65 184 66
rect 185 65 186 66
rect 20 140 21 141
rect 22 140 23 141
rect 23 140 24 141
rect 25 140 26 141
rect 20 141 26 145
rect 20 145 21 146
rect 22 145 23 146
rect 23 145 24 146
rect 25 145 26 146
rect 40 120 41 121
rect 42 120 43 121
rect 43 120 44 121
rect 45 120 46 121
rect 40 121 46 125
rect 40 125 41 126
rect 42 125 43 126
rect 43 125 44 126
rect 45 125 46 126
rect 380 260 381 261
rect 382 260 383 261
rect 383 260 384 261
rect 385 260 386 261
rect 380 261 386 265
rect 380 265 381 266
rect 382 265 383 266
rect 383 265 384 266
rect 385 265 386 266
rect 220 420 221 421
rect 222 420 223 421
rect 223 420 224 421
rect 225 420 226 421
rect 220 421 226 425
rect 220 425 221 426
rect 222 425 223 426
rect 223 425 224 426
rect 225 425 226 426
rect 300 120 301 121
rect 302 120 303 121
rect 303 120 304 121
rect 305 120 306 121
rect 300 121 306 125
rect 300 125 301 126
rect 302 125 303 126
rect 303 125 304 126
rect 305 125 306 126
rect 220 40 221 41
rect 222 40 223 41
rect 223 40 224 41
rect 225 40 226 41
rect 220 41 226 45
rect 220 45 221 46
rect 222 45 223 46
rect 223 45 224 46
rect 225 45 226 46
rect 200 160 201 161
rect 202 160 203 161
rect 203 160 204 161
rect 205 160 206 161
rect 200 161 206 165
rect 200 165 201 166
rect 202 165 203 166
rect 203 165 204 166
rect 205 165 206 166
rect 20 120 21 121
rect 22 120 23 121
rect 23 120 24 121
rect 25 120 26 121
rect 20 121 26 125
rect 20 125 21 126
rect 22 125 23 126
rect 23 125 24 126
rect 25 125 26 126
rect 160 240 161 241
rect 162 240 163 241
rect 163 240 164 241
rect 165 240 166 241
rect 160 241 166 245
rect 160 245 161 246
rect 162 245 163 246
rect 163 245 164 246
rect 165 245 166 246
rect 320 420 321 421
rect 322 420 323 421
rect 323 420 324 421
rect 325 420 326 421
rect 320 421 326 425
rect 320 425 321 426
rect 322 425 323 426
rect 323 425 324 426
rect 325 425 326 426
rect 220 20 221 21
rect 222 20 223 21
rect 223 20 224 21
rect 225 20 226 21
rect 220 21 226 25
rect 220 25 221 26
rect 222 25 223 26
rect 223 25 224 26
rect 225 25 226 26
rect 220 80 221 81
rect 222 80 223 81
rect 223 80 224 81
rect 225 80 226 81
rect 220 81 226 85
rect 220 85 221 86
rect 222 85 223 86
rect 223 85 224 86
rect 225 85 226 86
rect 320 160 321 161
rect 322 160 323 161
rect 323 160 324 161
rect 325 160 326 161
rect 320 161 326 165
rect 320 165 321 166
rect 322 165 323 166
rect 323 165 324 166
rect 325 165 326 166
rect 140 200 141 201
rect 142 200 143 201
rect 143 200 144 201
rect 145 200 146 201
rect 140 201 146 205
rect 140 205 141 206
rect 142 205 143 206
rect 143 205 144 206
rect 145 205 146 206
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect 400 220 401 221
rect 402 220 403 221
rect 403 220 404 221
rect 405 220 406 221
rect 400 221 406 225
rect 400 225 401 226
rect 402 225 403 226
rect 403 225 404 226
rect 405 225 406 226
rect 180 280 181 281
rect 182 280 183 281
rect 183 280 184 281
rect 185 280 186 281
rect 180 281 186 285
rect 180 285 181 286
rect 182 285 183 286
rect 183 285 184 286
rect 185 285 186 286
rect 200 300 201 301
rect 202 300 203 301
rect 203 300 204 301
rect 205 300 206 301
rect 200 301 206 305
rect 200 305 201 306
rect 202 305 203 306
rect 203 305 204 306
rect 205 305 206 306
rect 300 440 301 441
rect 302 440 303 441
rect 303 440 304 441
rect 305 440 306 441
rect 300 441 306 445
rect 300 445 301 446
rect 302 445 303 446
rect 303 445 304 446
rect 305 445 306 446
rect 100 260 101 261
rect 102 260 103 261
rect 103 260 104 261
rect 105 260 106 261
rect 100 261 106 265
rect 100 265 101 266
rect 102 265 103 266
rect 103 265 104 266
rect 105 265 106 266
rect 340 80 341 81
rect 342 80 343 81
rect 343 80 344 81
rect 345 80 346 81
rect 340 81 346 85
rect 340 85 341 86
rect 342 85 343 86
rect 343 85 344 86
rect 345 85 346 86
rect 160 0 161 1
rect 162 0 163 1
rect 163 0 164 1
rect 165 0 166 1
rect 160 1 166 5
rect 160 5 161 6
rect 162 5 163 6
rect 163 5 164 6
rect 165 5 166 6
rect 40 300 41 301
rect 42 300 43 301
rect 43 300 44 301
rect 45 300 46 301
rect 40 301 46 305
rect 40 305 41 306
rect 42 305 43 306
rect 43 305 44 306
rect 45 305 46 306
rect 140 260 141 261
rect 142 260 143 261
rect 143 260 144 261
rect 145 260 146 261
rect 140 261 146 265
rect 140 265 141 266
rect 142 265 143 266
rect 143 265 144 266
rect 145 265 146 266
rect 240 20 241 21
rect 242 20 243 21
rect 243 20 244 21
rect 245 20 246 21
rect 240 21 246 25
rect 240 25 241 26
rect 242 25 243 26
rect 243 25 244 26
rect 245 25 246 26
rect 140 380 141 381
rect 142 380 143 381
rect 143 380 144 381
rect 145 380 146 381
rect 140 381 146 385
rect 140 385 141 386
rect 142 385 143 386
rect 143 385 144 386
rect 145 385 146 386
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect 240 80 241 81
rect 242 80 243 81
rect 243 80 244 81
rect 245 80 246 81
rect 240 81 246 85
rect 240 85 241 86
rect 242 85 243 86
rect 243 85 244 86
rect 245 85 246 86
rect 40 260 41 261
rect 42 260 43 261
rect 43 260 44 261
rect 45 260 46 261
rect 40 261 46 265
rect 40 265 41 266
rect 42 265 43 266
rect 43 265 44 266
rect 45 265 46 266
rect 120 100 121 101
rect 122 100 123 101
rect 123 100 124 101
rect 125 100 126 101
rect 120 101 126 105
rect 120 105 121 106
rect 122 105 123 106
rect 123 105 124 106
rect 125 105 126 106
rect 320 80 321 81
rect 322 80 323 81
rect 323 80 324 81
rect 325 80 326 81
rect 320 81 326 85
rect 320 85 321 86
rect 322 85 323 86
rect 323 85 324 86
rect 325 85 326 86
rect 320 180 321 181
rect 322 180 323 181
rect 323 180 324 181
rect 325 180 326 181
rect 320 181 326 185
rect 320 185 321 186
rect 322 185 323 186
rect 323 185 324 186
rect 325 185 326 186
rect 280 340 281 341
rect 282 340 283 341
rect 283 340 284 341
rect 285 340 286 341
rect 280 341 286 345
rect 280 345 281 346
rect 282 345 283 346
rect 283 345 284 346
rect 285 345 286 346
rect 220 400 221 401
rect 222 400 223 401
rect 223 400 224 401
rect 225 400 226 401
rect 220 401 226 405
rect 220 405 221 406
rect 222 405 223 406
rect 223 405 224 406
rect 225 405 226 406
rect 100 180 101 181
rect 102 180 103 181
rect 103 180 104 181
rect 105 180 106 181
rect 100 181 106 185
rect 100 185 101 186
rect 102 185 103 186
rect 103 185 104 186
rect 105 185 106 186
rect 180 400 181 401
rect 182 400 183 401
rect 183 400 184 401
rect 185 400 186 401
rect 180 401 186 405
rect 180 405 181 406
rect 182 405 183 406
rect 183 405 184 406
rect 185 405 186 406
rect 180 440 181 441
rect 182 440 183 441
rect 183 440 184 441
rect 185 440 186 441
rect 180 441 186 445
rect 180 445 181 446
rect 182 445 183 446
rect 183 445 184 446
rect 185 445 186 446
rect 220 380 221 381
rect 222 380 223 381
rect 223 380 224 381
rect 225 380 226 381
rect 220 381 226 385
rect 220 385 221 386
rect 222 385 223 386
rect 223 385 224 386
rect 225 385 226 386
rect 400 120 401 121
rect 402 120 403 121
rect 403 120 404 121
rect 405 120 406 121
rect 400 121 406 125
rect 400 125 401 126
rect 402 125 403 126
rect 403 125 404 126
rect 405 125 406 126
rect 380 200 381 201
rect 382 200 383 201
rect 383 200 384 201
rect 385 200 386 201
rect 380 201 386 205
rect 380 205 381 206
rect 382 205 383 206
rect 383 205 384 206
rect 385 205 386 206
rect 260 180 261 181
rect 262 180 263 181
rect 263 180 264 181
rect 265 180 266 181
rect 260 181 266 185
rect 260 185 261 186
rect 262 185 263 186
rect 263 185 264 186
rect 265 185 266 186
rect 340 120 341 121
rect 342 120 343 121
rect 343 120 344 121
rect 345 120 346 121
rect 340 121 346 125
rect 340 125 341 126
rect 342 125 343 126
rect 343 125 344 126
rect 345 125 346 126
rect 160 400 161 401
rect 162 400 163 401
rect 163 400 164 401
rect 165 400 166 401
rect 160 401 166 405
rect 160 405 161 406
rect 162 405 163 406
rect 163 405 164 406
rect 165 405 166 406
rect 0 100 1 101
rect 2 100 3 101
rect 3 100 4 101
rect 5 100 6 101
rect 0 101 6 105
rect 0 105 1 106
rect 2 105 3 106
rect 3 105 4 106
rect 5 105 6 106
rect 80 60 81 61
rect 82 60 83 61
rect 83 60 84 61
rect 85 60 86 61
rect 80 61 86 65
rect 80 65 81 66
rect 82 65 83 66
rect 83 65 84 66
rect 85 65 86 66
rect 0 160 1 161
rect 2 160 3 161
rect 3 160 4 161
rect 5 160 6 161
rect 0 161 6 165
rect 0 165 1 166
rect 2 165 3 166
rect 3 165 4 166
rect 5 165 6 166
rect 280 460 281 461
rect 282 460 283 461
rect 283 460 284 461
rect 285 460 286 461
rect 280 461 286 465
rect 280 465 281 466
rect 282 465 283 466
rect 283 465 284 466
rect 285 465 286 466
rect 160 140 161 141
rect 162 140 163 141
rect 163 140 164 141
rect 165 140 166 141
rect 160 141 166 145
rect 160 145 161 146
rect 162 145 163 146
rect 163 145 164 146
rect 165 145 166 146
rect 180 300 181 301
rect 182 300 183 301
rect 183 300 184 301
rect 185 300 186 301
rect 180 301 186 305
rect 180 305 181 306
rect 182 305 183 306
rect 183 305 184 306
rect 185 305 186 306
rect 420 180 421 181
rect 422 180 423 181
rect 423 180 424 181
rect 425 180 426 181
rect 420 181 426 185
rect 420 185 421 186
rect 422 185 423 186
rect 423 185 424 186
rect 425 185 426 186
rect 140 340 141 341
rect 142 340 143 341
rect 143 340 144 341
rect 145 340 146 341
rect 140 341 146 345
rect 140 345 141 346
rect 142 345 143 346
rect 143 345 144 346
rect 145 345 146 346
rect 360 320 361 321
rect 362 320 363 321
rect 363 320 364 321
rect 365 320 366 321
rect 360 321 366 325
rect 360 325 361 326
rect 362 325 363 326
rect 363 325 364 326
rect 365 325 366 326
rect 280 120 281 121
rect 282 120 283 121
rect 283 120 284 121
rect 285 120 286 121
rect 280 121 286 125
rect 280 125 281 126
rect 282 125 283 126
rect 283 125 284 126
rect 285 125 286 126
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect 140 360 141 361
rect 142 360 143 361
rect 143 360 144 361
rect 145 360 146 361
rect 140 361 146 365
rect 140 365 141 366
rect 142 365 143 366
rect 143 365 144 366
rect 145 365 146 366
rect 180 100 181 101
rect 182 100 183 101
rect 183 100 184 101
rect 185 100 186 101
rect 180 101 186 105
rect 180 105 181 106
rect 182 105 183 106
rect 183 105 184 106
rect 185 105 186 106
rect 100 40 101 41
rect 102 40 103 41
rect 103 40 104 41
rect 105 40 106 41
rect 100 41 106 45
rect 100 45 101 46
rect 102 45 103 46
rect 103 45 104 46
rect 105 45 106 46
rect 100 60 101 61
rect 102 60 103 61
rect 103 60 104 61
rect 105 60 106 61
rect 100 61 106 65
rect 100 65 101 66
rect 102 65 103 66
rect 103 65 104 66
rect 105 65 106 66
rect 260 260 261 261
rect 262 260 263 261
rect 263 260 264 261
rect 265 260 266 261
rect 260 261 266 265
rect 260 265 261 266
rect 262 265 263 266
rect 263 265 264 266
rect 265 265 266 266
rect 240 380 241 381
rect 242 380 243 381
rect 243 380 244 381
rect 245 380 246 381
rect 240 381 246 385
rect 240 385 241 386
rect 242 385 243 386
rect 243 385 244 386
rect 245 385 246 386
rect 20 240 21 241
rect 22 240 23 241
rect 23 240 24 241
rect 25 240 26 241
rect 20 241 26 245
rect 20 245 21 246
rect 22 245 23 246
rect 23 245 24 246
rect 25 245 26 246
rect 60 120 61 121
rect 62 120 63 121
rect 63 120 64 121
rect 65 120 66 121
rect 60 121 66 125
rect 60 125 61 126
rect 62 125 63 126
rect 63 125 64 126
rect 65 125 66 126
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect 180 260 181 261
rect 182 260 183 261
rect 183 260 184 261
rect 185 260 186 261
rect 180 261 186 265
rect 180 265 181 266
rect 182 265 183 266
rect 183 265 184 266
rect 185 265 186 266
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect 220 320 221 321
rect 222 320 223 321
rect 223 320 224 321
rect 225 320 226 321
rect 220 321 226 325
rect 220 325 221 326
rect 222 325 223 326
rect 223 325 224 326
rect 225 325 226 326
rect 160 420 161 421
rect 162 420 163 421
rect 163 420 164 421
rect 165 420 166 421
rect 160 421 166 425
rect 160 425 161 426
rect 162 425 163 426
rect 163 425 164 426
rect 165 425 166 426
rect 320 440 321 441
rect 322 440 323 441
rect 323 440 324 441
rect 325 440 326 441
rect 320 441 326 445
rect 320 445 321 446
rect 322 445 323 446
rect 323 445 324 446
rect 325 445 326 446
rect 100 120 101 121
rect 102 120 103 121
rect 103 120 104 121
rect 105 120 106 121
rect 100 121 106 125
rect 100 125 101 126
rect 102 125 103 126
rect 103 125 104 126
rect 105 125 106 126
rect 280 220 281 221
rect 282 220 283 221
rect 283 220 284 221
rect 285 220 286 221
rect 280 221 286 225
rect 280 225 281 226
rect 282 225 283 226
rect 283 225 284 226
rect 285 225 286 226
rect 140 420 141 421
rect 142 420 143 421
rect 143 420 144 421
rect 145 420 146 421
rect 140 421 146 425
rect 140 425 141 426
rect 142 425 143 426
rect 143 425 144 426
rect 145 425 146 426
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect 260 100 261 101
rect 262 100 263 101
rect 263 100 264 101
rect 265 100 266 101
rect 260 101 266 105
rect 260 105 261 106
rect 262 105 263 106
rect 263 105 264 106
rect 265 105 266 106
rect 240 100 241 101
rect 242 100 243 101
rect 243 100 244 101
rect 245 100 246 101
rect 240 101 246 105
rect 240 105 241 106
rect 242 105 243 106
rect 243 105 244 106
rect 245 105 246 106
rect 80 240 81 241
rect 82 240 83 241
rect 83 240 84 241
rect 85 240 86 241
rect 80 241 86 245
rect 80 245 81 246
rect 82 245 83 246
rect 83 245 84 246
rect 85 245 86 246
rect 340 360 341 361
rect 342 360 343 361
rect 343 360 344 361
rect 345 360 346 361
rect 340 361 346 365
rect 340 365 341 366
rect 342 365 343 366
rect 343 365 344 366
rect 345 365 346 366
rect 240 340 241 341
rect 242 340 243 341
rect 243 340 244 341
rect 245 340 246 341
rect 240 341 246 345
rect 240 345 241 346
rect 242 345 243 346
rect 243 345 244 346
rect 245 345 246 346
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect 240 220 241 221
rect 242 220 243 221
rect 243 220 244 221
rect 245 220 246 221
rect 240 221 246 225
rect 240 225 241 226
rect 242 225 243 226
rect 243 225 244 226
rect 245 225 246 226
rect 300 140 301 141
rect 302 140 303 141
rect 303 140 304 141
rect 305 140 306 141
rect 300 141 306 145
rect 300 145 301 146
rect 302 145 303 146
rect 303 145 304 146
rect 305 145 306 146
rect 240 60 241 61
rect 242 60 243 61
rect 243 60 244 61
rect 245 60 246 61
rect 240 61 246 65
rect 240 65 241 66
rect 242 65 243 66
rect 243 65 244 66
rect 245 65 246 66
rect 20 200 21 201
rect 22 200 23 201
rect 23 200 24 201
rect 25 200 26 201
rect 20 201 26 205
rect 20 205 21 206
rect 22 205 23 206
rect 23 205 24 206
rect 25 205 26 206
rect 140 140 141 141
rect 142 140 143 141
rect 143 140 144 141
rect 145 140 146 141
rect 140 141 146 145
rect 140 145 141 146
rect 142 145 143 146
rect 143 145 144 146
rect 145 145 146 146
rect 260 20 261 21
rect 262 20 263 21
rect 263 20 264 21
rect 265 20 266 21
rect 260 21 266 25
rect 260 25 261 26
rect 262 25 263 26
rect 263 25 264 26
rect 265 25 266 26
rect 360 180 361 181
rect 362 180 363 181
rect 363 180 364 181
rect 365 180 366 181
rect 360 181 366 185
rect 360 185 361 186
rect 362 185 363 186
rect 363 185 364 186
rect 365 185 366 186
rect 300 420 301 421
rect 302 420 303 421
rect 303 420 304 421
rect 305 420 306 421
rect 300 421 306 425
rect 300 425 301 426
rect 302 425 303 426
rect 303 425 304 426
rect 305 425 306 426
rect 200 360 201 361
rect 202 360 203 361
rect 203 360 204 361
rect 205 360 206 361
rect 200 361 206 365
rect 200 365 201 366
rect 202 365 203 366
rect 203 365 204 366
rect 205 365 206 366
rect 100 200 101 201
rect 102 200 103 201
rect 103 200 104 201
rect 105 200 106 201
rect 100 201 106 205
rect 100 205 101 206
rect 102 205 103 206
rect 103 205 104 206
rect 105 205 106 206
rect 160 380 161 381
rect 162 380 163 381
rect 163 380 164 381
rect 165 380 166 381
rect 160 381 166 385
rect 160 385 161 386
rect 162 385 163 386
rect 163 385 164 386
rect 165 385 166 386
rect 260 320 261 321
rect 262 320 263 321
rect 263 320 264 321
rect 265 320 266 321
rect 260 321 266 325
rect 260 325 261 326
rect 262 325 263 326
rect 263 325 264 326
rect 265 325 266 326
rect 380 240 381 241
rect 382 240 383 241
rect 383 240 384 241
rect 385 240 386 241
rect 380 241 386 245
rect 380 245 381 246
rect 382 245 383 246
rect 383 245 384 246
rect 385 245 386 246
rect 40 280 41 281
rect 42 280 43 281
rect 43 280 44 281
rect 45 280 46 281
rect 40 281 46 285
rect 40 285 41 286
rect 42 285 43 286
rect 43 285 44 286
rect 45 285 46 286
rect 300 60 301 61
rect 302 60 303 61
rect 303 60 304 61
rect 305 60 306 61
rect 300 61 306 65
rect 300 65 301 66
rect 302 65 303 66
rect 303 65 304 66
rect 305 65 306 66
rect 100 280 101 281
rect 102 280 103 281
rect 103 280 104 281
rect 105 280 106 281
rect 100 281 106 285
rect 100 285 101 286
rect 102 285 103 286
rect 103 285 104 286
rect 105 285 106 286
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect 80 260 81 261
rect 82 260 83 261
rect 83 260 84 261
rect 85 260 86 261
rect 80 261 86 265
rect 80 265 81 266
rect 82 265 83 266
rect 83 265 84 266
rect 85 265 86 266
rect 380 180 381 181
rect 382 180 383 181
rect 383 180 384 181
rect 385 180 386 181
rect 380 181 386 185
rect 380 185 381 186
rect 382 185 383 186
rect 383 185 384 186
rect 385 185 386 186
rect 380 360 381 361
rect 382 360 383 361
rect 383 360 384 361
rect 385 360 386 361
rect 380 361 386 365
rect 380 365 381 366
rect 382 365 383 366
rect 383 365 384 366
rect 385 365 386 366
rect 140 300 141 301
rect 142 300 143 301
rect 143 300 144 301
rect 145 300 146 301
rect 140 301 146 305
rect 140 305 141 306
rect 142 305 143 306
rect 143 305 144 306
rect 145 305 146 306
rect 340 260 341 261
rect 342 260 343 261
rect 343 260 344 261
rect 345 260 346 261
rect 340 261 346 265
rect 340 265 341 266
rect 342 265 343 266
rect 343 265 344 266
rect 345 265 346 266
rect 100 360 101 361
rect 102 360 103 361
rect 103 360 104 361
rect 105 360 106 361
rect 100 361 106 365
rect 100 365 101 366
rect 102 365 103 366
rect 103 365 104 366
rect 105 365 106 366
rect 140 220 141 221
rect 142 220 143 221
rect 143 220 144 221
rect 145 220 146 221
rect 140 221 146 225
rect 140 225 141 226
rect 142 225 143 226
rect 143 225 144 226
rect 145 225 146 226
rect 240 420 241 421
rect 242 420 243 421
rect 243 420 244 421
rect 245 420 246 421
rect 240 421 246 425
rect 240 425 241 426
rect 242 425 243 426
rect 243 425 244 426
rect 245 425 246 426
<< polysilicon >>
rect 121 319 122 321
rect 124 319 125 321
rect 121 325 122 327
rect 124 325 125 327
rect 361 239 362 241
rect 364 239 365 241
rect 361 245 362 247
rect 364 245 365 247
rect 141 319 142 321
rect 144 319 145 321
rect 141 325 142 327
rect 144 325 145 327
rect 261 359 262 361
rect 264 359 265 361
rect 261 365 262 367
rect 264 365 265 367
rect 181 379 182 381
rect 184 379 185 381
rect 181 385 182 387
rect 184 385 185 387
rect 321 239 322 241
rect 324 239 325 241
rect 321 245 322 247
rect 324 245 325 247
rect 81 399 82 401
rect 84 399 85 401
rect 81 405 82 407
rect 84 405 85 407
rect 81 299 82 301
rect 84 299 85 301
rect 81 305 82 307
rect 84 305 85 307
rect 361 159 362 161
rect 364 159 365 161
rect 361 165 362 167
rect 364 165 365 167
rect 321 199 322 201
rect 324 199 325 201
rect 321 205 322 207
rect 324 205 325 207
rect 321 319 322 321
rect 324 319 325 321
rect 321 325 322 327
rect 324 325 325 327
rect 381 159 382 161
rect 384 159 385 161
rect 381 165 382 167
rect 384 165 385 167
rect 281 399 282 401
rect 284 399 285 401
rect 281 405 282 407
rect 284 405 285 407
rect 1 139 2 141
rect 4 139 5 141
rect 1 145 2 147
rect 4 145 5 147
rect 101 339 102 341
rect 104 339 105 341
rect 101 345 102 347
rect 104 345 105 347
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect 81 279 82 281
rect 84 279 85 281
rect 81 285 82 287
rect 84 285 85 287
rect 121 359 122 361
rect 124 359 125 361
rect 121 365 122 367
rect 124 365 125 367
rect 81 159 82 161
rect 84 159 85 161
rect 81 165 82 167
rect 84 165 85 167
rect 321 219 322 221
rect 324 219 325 221
rect 321 225 322 227
rect 324 225 325 227
rect 261 439 262 441
rect 264 439 265 441
rect 261 445 262 447
rect 264 445 265 447
rect 201 279 202 281
rect 204 279 205 281
rect 201 285 202 287
rect 204 285 205 287
rect 361 259 362 261
rect 364 259 365 261
rect 361 265 362 267
rect 364 265 365 267
rect 401 239 402 241
rect 404 239 405 241
rect 401 245 402 247
rect 404 245 405 247
rect 81 119 82 121
rect 84 119 85 121
rect 81 125 82 127
rect 84 125 85 127
rect 321 399 322 401
rect 324 399 325 401
rect 321 405 322 407
rect 324 405 325 407
rect 261 299 262 301
rect 264 299 265 301
rect 261 305 262 307
rect 264 305 265 307
rect 161 299 162 301
rect 164 299 165 301
rect 161 305 162 307
rect 164 305 165 307
rect 261 39 262 41
rect 264 39 265 41
rect 261 45 262 47
rect 264 45 265 47
rect 241 259 242 261
rect 244 259 245 261
rect 241 265 242 267
rect 244 265 245 267
rect 181 119 182 121
rect 184 119 185 121
rect 181 125 182 127
rect 184 125 185 127
rect 41 139 42 141
rect 44 139 45 141
rect 41 145 42 147
rect 44 145 45 147
rect 401 259 402 261
rect 404 259 405 261
rect 401 265 402 267
rect 404 265 405 267
rect 241 299 242 301
rect 244 299 245 301
rect 241 305 242 307
rect 244 305 245 307
rect 161 179 162 181
rect 164 179 165 181
rect 161 185 162 187
rect 164 185 165 187
rect 261 339 262 341
rect 264 339 265 341
rect 261 345 262 347
rect 264 345 265 347
rect 121 239 122 241
rect 124 239 125 241
rect 121 245 122 247
rect 124 245 125 247
rect 401 159 402 161
rect 404 159 405 161
rect 401 165 402 167
rect 404 165 405 167
rect 41 159 42 161
rect 44 159 45 161
rect 41 165 42 167
rect 44 165 45 167
rect 281 379 282 381
rect 284 379 285 381
rect 281 385 282 387
rect 284 385 285 387
rect 141 399 142 401
rect 144 399 145 401
rect 141 405 142 407
rect 144 405 145 407
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect 281 99 282 101
rect 284 99 285 101
rect 281 105 282 107
rect 284 105 285 107
rect 101 79 102 81
rect 104 79 105 81
rect 101 85 102 87
rect 104 85 105 87
rect 401 199 402 201
rect 404 199 405 201
rect 401 205 402 207
rect 404 205 405 207
rect 281 299 282 301
rect 284 299 285 301
rect 281 305 282 307
rect 284 305 285 307
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect 281 439 282 441
rect 284 439 285 441
rect 281 445 282 447
rect 284 445 285 447
rect 161 339 162 341
rect 164 339 165 341
rect 161 345 162 347
rect 164 345 165 347
rect 101 99 102 101
rect 104 99 105 101
rect 101 105 102 107
rect 104 105 105 107
rect 201 219 202 221
rect 204 219 205 221
rect 201 225 202 227
rect 204 225 205 227
rect 101 319 102 321
rect 104 319 105 321
rect 101 325 102 327
rect 104 325 105 327
rect 161 259 162 261
rect 164 259 165 261
rect 161 265 162 267
rect 164 265 165 267
rect 121 199 122 201
rect 124 199 125 201
rect 121 205 122 207
rect 124 205 125 207
rect 281 59 282 61
rect 284 59 285 61
rect 281 65 282 67
rect 284 65 285 67
rect 81 319 82 321
rect 84 319 85 321
rect 81 325 82 327
rect 84 325 85 327
rect 361 359 362 361
rect 364 359 365 361
rect 361 365 362 367
rect 364 365 365 367
rect 201 119 202 121
rect 204 119 205 121
rect 201 125 202 127
rect 204 125 205 127
rect 241 279 242 281
rect 244 279 245 281
rect 241 285 242 287
rect 244 285 245 287
rect 261 219 262 221
rect 264 219 265 221
rect 261 225 262 227
rect 264 225 265 227
rect 221 199 222 201
rect 224 199 225 201
rect 221 205 222 207
rect 224 205 225 207
rect 261 399 262 401
rect 264 399 265 401
rect 261 405 262 407
rect 264 405 265 407
rect 141 239 142 241
rect 144 239 145 241
rect 141 245 142 247
rect 144 245 145 247
rect 241 159 242 161
rect 244 159 245 161
rect 241 165 242 167
rect 244 165 245 167
rect 101 239 102 241
rect 104 239 105 241
rect 101 245 102 247
rect 104 245 105 247
rect 161 319 162 321
rect 164 319 165 321
rect 161 325 162 327
rect 164 325 165 327
rect 161 159 162 161
rect 164 159 165 161
rect 161 165 162 167
rect 164 165 165 167
rect 81 359 82 361
rect 84 359 85 361
rect 81 365 82 367
rect 84 365 85 367
rect 41 99 42 101
rect 44 99 45 101
rect 41 105 42 107
rect 44 105 45 107
rect 201 439 202 441
rect 204 439 205 441
rect 201 445 202 447
rect 204 445 205 447
rect 61 199 62 201
rect 64 199 65 201
rect 61 205 62 207
rect 64 205 65 207
rect 1 179 2 181
rect 4 179 5 181
rect 1 185 2 187
rect 4 185 5 187
rect 181 199 182 201
rect 184 199 185 201
rect 181 205 182 207
rect 184 205 185 207
rect 301 399 302 401
rect 304 399 305 401
rect 301 405 302 407
rect 304 405 305 407
rect 301 159 302 161
rect 304 159 305 161
rect 301 165 302 167
rect 304 165 305 167
rect 1 219 2 221
rect 4 219 5 221
rect 1 225 2 227
rect 4 225 5 227
rect 381 139 382 141
rect 384 139 385 141
rect 381 145 382 147
rect 384 145 385 147
rect 81 39 82 41
rect 84 39 85 41
rect 81 45 82 47
rect 84 45 85 47
rect 121 339 122 341
rect 124 339 125 341
rect 121 345 122 347
rect 124 345 125 347
rect 61 299 62 301
rect 64 299 65 301
rect 61 305 62 307
rect 64 305 65 307
rect 241 -1 242 1
rect 244 -1 245 1
rect 241 5 242 7
rect 244 5 245 7
rect 281 239 282 241
rect 284 239 285 241
rect 281 245 282 247
rect 284 245 285 247
rect 41 319 42 321
rect 44 319 45 321
rect 41 325 42 327
rect 44 325 45 327
rect 201 99 202 101
rect 204 99 205 101
rect 201 105 202 107
rect 204 105 205 107
rect 301 99 302 101
rect 304 99 305 101
rect 301 105 302 107
rect 304 105 305 107
rect 321 299 322 301
rect 324 299 325 301
rect 321 305 322 307
rect 324 305 325 307
rect 1 119 2 121
rect 4 119 5 121
rect 1 125 2 127
rect 4 125 5 127
rect 421 239 422 241
rect 424 239 425 241
rect 421 245 422 247
rect 424 245 425 247
rect 301 339 302 341
rect 304 339 305 341
rect 301 345 302 347
rect 304 345 305 347
rect 161 199 162 201
rect 164 199 165 201
rect 161 205 162 207
rect 164 205 165 207
rect 101 139 102 141
rect 104 139 105 141
rect 101 145 102 147
rect 104 145 105 147
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect 381 279 382 281
rect 384 279 385 281
rect 381 285 382 287
rect 384 285 385 287
rect 21 159 22 161
rect 24 159 25 161
rect 21 165 22 167
rect 24 165 25 167
rect 121 179 122 181
rect 124 179 125 181
rect 121 185 122 187
rect 124 185 125 187
rect 121 119 122 121
rect 124 119 125 121
rect 121 125 122 127
rect 124 125 125 127
rect 421 199 422 201
rect 424 199 425 201
rect 421 205 422 207
rect 424 205 425 207
rect 221 239 222 241
rect 224 239 225 241
rect 221 245 222 247
rect 224 245 225 247
rect 241 239 242 241
rect 244 239 245 241
rect 241 245 242 247
rect 244 245 245 247
rect 421 219 422 221
rect 424 219 425 221
rect 421 225 422 227
rect 424 225 425 227
rect 181 419 182 421
rect 184 419 185 421
rect 181 425 182 427
rect 184 425 185 427
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect 341 399 342 401
rect 344 399 345 401
rect 341 405 342 407
rect 344 405 345 407
rect 81 219 82 221
rect 84 219 85 221
rect 81 225 82 227
rect 84 225 85 227
rect 41 239 42 241
rect 44 239 45 241
rect 41 245 42 247
rect 44 245 45 247
rect 181 359 182 361
rect 184 359 185 361
rect 181 365 182 367
rect 184 365 185 367
rect 341 219 342 221
rect 344 219 345 221
rect 341 225 342 227
rect 344 225 345 227
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect 281 -1 282 1
rect 284 -1 285 1
rect 281 5 282 7
rect 284 5 285 7
rect 261 159 262 161
rect 264 159 265 161
rect 261 165 262 167
rect 264 165 265 167
rect 281 319 282 321
rect 284 319 285 321
rect 281 325 282 327
rect 284 325 285 327
rect 121 219 122 221
rect 124 219 125 221
rect 121 225 122 227
rect 124 225 125 227
rect 61 159 62 161
rect 64 159 65 161
rect 61 165 62 167
rect 64 165 65 167
rect 261 119 262 121
rect 264 119 265 121
rect 261 125 262 127
rect 264 125 265 127
rect 161 99 162 101
rect 164 99 165 101
rect 161 105 162 107
rect 164 105 165 107
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect 361 219 362 221
rect 364 219 365 221
rect 361 225 362 227
rect 364 225 365 227
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect 101 399 102 401
rect 104 399 105 401
rect 101 405 102 407
rect 104 405 105 407
rect 421 119 422 121
rect 424 119 425 121
rect 421 125 422 127
rect 424 125 425 127
rect 21 179 22 181
rect 24 179 25 181
rect 21 185 22 187
rect 24 185 25 187
rect 201 59 202 61
rect 204 59 205 61
rect 201 65 202 67
rect 204 65 205 67
rect 81 79 82 81
rect 84 79 85 81
rect 81 85 82 87
rect 84 85 85 87
rect 241 399 242 401
rect 244 399 245 401
rect 241 405 242 407
rect 244 405 245 407
rect 61 239 62 241
rect 64 239 65 241
rect 61 245 62 247
rect 64 245 65 247
rect 141 159 142 161
rect 144 159 145 161
rect 141 165 142 167
rect 144 165 145 167
rect 301 319 302 321
rect 304 319 305 321
rect 301 325 302 327
rect 304 325 305 327
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect 201 19 202 21
rect 204 19 205 21
rect 201 25 202 27
rect 204 25 205 27
rect 281 19 282 21
rect 284 19 285 21
rect 281 25 282 27
rect 284 25 285 27
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect 181 319 182 321
rect 184 319 185 321
rect 181 325 182 327
rect 184 325 185 327
rect 221 139 222 141
rect 224 139 225 141
rect 221 145 222 147
rect 224 145 225 147
rect 321 59 322 61
rect 324 59 325 61
rect 321 65 322 67
rect 324 65 325 67
rect 21 219 22 221
rect 24 219 25 221
rect 21 225 22 227
rect 24 225 25 227
rect 281 259 282 261
rect 284 259 285 261
rect 281 265 282 267
rect 284 265 285 267
rect 141 279 142 281
rect 144 279 145 281
rect 141 285 142 287
rect 144 285 145 287
rect 301 279 302 281
rect 304 279 305 281
rect 301 285 302 287
rect 304 285 305 287
rect 401 179 402 181
rect 404 179 405 181
rect 401 185 402 187
rect 404 185 405 187
rect 141 119 142 121
rect 144 119 145 121
rect 141 125 142 127
rect 144 125 145 127
rect 121 139 122 141
rect 124 139 125 141
rect 121 145 122 147
rect 124 145 125 147
rect 261 199 262 201
rect 264 199 265 201
rect 261 205 262 207
rect 264 205 265 207
rect 161 219 162 221
rect 164 219 165 221
rect 161 225 162 227
rect 164 225 165 227
rect 261 459 262 461
rect 264 459 265 461
rect 261 465 262 467
rect 264 465 265 467
rect 121 59 122 61
rect 124 59 125 61
rect 121 65 122 67
rect 124 65 125 67
rect 301 359 302 361
rect 304 359 305 361
rect 301 365 302 367
rect 304 365 305 367
rect 201 139 202 141
rect 204 139 205 141
rect 201 145 202 147
rect 204 145 205 147
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect 101 159 102 161
rect 104 159 105 161
rect 101 165 102 167
rect 104 165 105 167
rect 241 39 242 41
rect 244 39 245 41
rect 241 45 242 47
rect 244 45 245 47
rect 221 299 222 301
rect 224 299 225 301
rect 221 305 222 307
rect 224 305 225 307
rect 201 79 202 81
rect 204 79 205 81
rect 201 85 202 87
rect 204 85 205 87
rect 201 39 202 41
rect 204 39 205 41
rect 201 45 202 47
rect 204 45 205 47
rect 321 359 322 361
rect 324 359 325 361
rect 321 365 322 367
rect 324 365 325 367
rect 341 279 342 281
rect 344 279 345 281
rect 341 285 342 287
rect 344 285 345 287
rect 361 99 362 101
rect 364 99 365 101
rect 361 105 362 107
rect 364 105 365 107
rect 81 139 82 141
rect 84 139 85 141
rect 81 145 82 147
rect 84 145 85 147
rect 61 79 62 81
rect 64 79 65 81
rect 61 85 62 87
rect 64 85 65 87
rect 121 279 122 281
rect 124 279 125 281
rect 121 285 122 287
rect 124 285 125 287
rect 261 239 262 241
rect 264 239 265 241
rect 261 245 262 247
rect 264 245 265 247
rect 321 379 322 381
rect 324 379 325 381
rect 321 385 322 387
rect 324 385 325 387
rect 161 359 162 361
rect 164 359 165 361
rect 161 365 162 367
rect 164 365 165 367
rect 221 99 222 101
rect 224 99 225 101
rect 221 105 222 107
rect 224 105 225 107
rect 181 79 182 81
rect 184 79 185 81
rect 181 85 182 87
rect 184 85 185 87
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect 241 319 242 321
rect 244 319 245 321
rect 241 325 242 327
rect 244 325 245 327
rect 301 299 302 301
rect 304 299 305 301
rect 301 305 302 307
rect 304 305 305 307
rect 201 319 202 321
rect 204 319 205 321
rect 201 325 202 327
rect 204 325 205 327
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect 61 319 62 321
rect 64 319 65 321
rect 61 325 62 327
rect 64 325 65 327
rect 221 159 222 161
rect 224 159 225 161
rect 221 165 222 167
rect 224 165 225 167
rect 81 379 82 381
rect 84 379 85 381
rect 81 385 82 387
rect 84 385 85 387
rect 261 379 262 381
rect 264 379 265 381
rect 261 385 262 387
rect 264 385 265 387
rect 341 339 342 341
rect 344 339 345 341
rect 341 345 342 347
rect 344 345 345 347
rect 281 159 282 161
rect 284 159 285 161
rect 281 165 282 167
rect 284 165 285 167
rect 21 279 22 281
rect 24 279 25 281
rect 21 285 22 287
rect 24 285 25 287
rect 361 279 362 281
rect 364 279 365 281
rect 361 285 362 287
rect 364 285 365 287
rect 41 219 42 221
rect 44 219 45 221
rect 41 225 42 227
rect 44 225 45 227
rect 141 59 142 61
rect 144 59 145 61
rect 141 65 142 67
rect 144 65 145 67
rect 181 159 182 161
rect 184 159 185 161
rect 181 165 182 167
rect 184 165 185 167
rect 361 379 362 381
rect 364 379 365 381
rect 361 385 362 387
rect 364 385 365 387
rect 81 179 82 181
rect 84 179 85 181
rect 81 185 82 187
rect 84 185 85 187
rect 221 259 222 261
rect 224 259 225 261
rect 221 265 222 267
rect 224 265 225 267
rect 341 139 342 141
rect 344 139 345 141
rect 341 145 342 147
rect 344 145 345 147
rect 141 39 142 41
rect 144 39 145 41
rect 141 45 142 47
rect 144 45 145 47
rect 101 379 102 381
rect 104 379 105 381
rect 101 385 102 387
rect 104 385 105 387
rect 341 199 342 201
rect 344 199 345 201
rect 341 205 342 207
rect 344 205 345 207
rect 321 279 322 281
rect 324 279 325 281
rect 321 285 322 287
rect 324 285 325 287
rect 201 259 202 261
rect 204 259 205 261
rect 201 265 202 267
rect 204 265 205 267
rect 201 399 202 401
rect 204 399 205 401
rect 201 405 202 407
rect 204 405 205 407
rect 81 99 82 101
rect 84 99 85 101
rect 81 105 82 107
rect 84 105 85 107
rect 61 99 62 101
rect 64 99 65 101
rect 61 105 62 107
rect 64 105 65 107
rect 141 79 142 81
rect 144 79 145 81
rect 141 85 142 87
rect 144 85 145 87
rect 281 139 282 141
rect 284 139 285 141
rect 281 145 282 147
rect 284 145 285 147
rect 301 179 302 181
rect 304 179 305 181
rect 301 185 302 187
rect 304 185 305 187
rect 341 299 342 301
rect 344 299 345 301
rect 341 305 342 307
rect 344 305 345 307
rect 401 299 402 301
rect 404 299 405 301
rect 401 305 402 307
rect 404 305 405 307
rect 221 359 222 361
rect 224 359 225 361
rect 221 365 222 367
rect 224 365 225 367
rect 181 219 182 221
rect 184 219 185 221
rect 181 225 182 227
rect 184 225 185 227
rect 161 59 162 61
rect 164 59 165 61
rect 161 65 162 67
rect 164 65 165 67
rect 41 179 42 181
rect 44 179 45 181
rect 41 185 42 187
rect 44 185 45 187
rect 61 279 62 281
rect 64 279 65 281
rect 61 285 62 287
rect 64 285 65 287
rect 181 179 182 181
rect 184 179 185 181
rect 181 185 182 187
rect 184 185 185 187
rect 161 119 162 121
rect 164 119 165 121
rect 161 125 162 127
rect 164 125 165 127
rect 381 319 382 321
rect 384 319 385 321
rect 381 325 382 327
rect 384 325 385 327
rect 241 199 242 201
rect 244 199 245 201
rect 241 205 242 207
rect 244 205 245 207
rect 81 339 82 341
rect 84 339 85 341
rect 81 345 82 347
rect 84 345 85 347
rect 361 299 362 301
rect 364 299 365 301
rect 361 305 362 307
rect 364 305 365 307
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect 301 379 302 381
rect 304 379 305 381
rect 301 385 302 387
rect 304 385 305 387
rect 321 259 322 261
rect 324 259 325 261
rect 321 265 322 267
rect 324 265 325 267
rect 341 239 342 241
rect 344 239 345 241
rect 341 245 342 247
rect 344 245 345 247
rect 121 159 122 161
rect 124 159 125 161
rect 121 165 122 167
rect 124 165 125 167
rect 281 179 282 181
rect 284 179 285 181
rect 281 185 282 187
rect 284 185 285 187
rect 221 339 222 341
rect 224 339 225 341
rect 221 345 222 347
rect 224 345 225 347
rect 101 219 102 221
rect 104 219 105 221
rect 101 225 102 227
rect 104 225 105 227
rect 181 139 182 141
rect 184 139 185 141
rect 181 145 182 147
rect 184 145 185 147
rect 361 339 362 341
rect 364 339 365 341
rect 361 345 362 347
rect 364 345 365 347
rect 61 219 62 221
rect 64 219 65 221
rect 61 225 62 227
rect 64 225 65 227
rect 281 279 282 281
rect 284 279 285 281
rect 281 285 282 287
rect 284 285 285 287
rect 321 99 322 101
rect 324 99 325 101
rect 321 105 322 107
rect 324 105 325 107
rect 381 219 382 221
rect 384 219 385 221
rect 381 225 382 227
rect 384 225 385 227
rect 121 79 122 81
rect 124 79 125 81
rect 121 85 122 87
rect 124 85 125 87
rect 321 139 322 141
rect 324 139 325 141
rect 321 145 322 147
rect 324 145 325 147
rect 1 259 2 261
rect 4 259 5 261
rect 1 265 2 267
rect 4 265 5 267
rect 321 39 322 41
rect 324 39 325 41
rect 321 45 322 47
rect 324 45 325 47
rect 221 219 222 221
rect 224 219 225 221
rect 221 225 222 227
rect 224 225 225 227
rect 101 299 102 301
rect 104 299 105 301
rect 101 305 102 307
rect 104 305 105 307
rect 281 79 282 81
rect 284 79 285 81
rect 281 85 282 87
rect 284 85 285 87
rect 181 19 182 21
rect 184 19 185 21
rect 181 25 182 27
rect 184 25 185 27
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect 221 59 222 61
rect 224 59 225 61
rect 221 65 222 67
rect 224 65 225 67
rect 201 199 202 201
rect 204 199 205 201
rect 201 205 202 207
rect 204 205 205 207
rect 261 139 262 141
rect 264 139 265 141
rect 261 145 262 147
rect 264 145 265 147
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect 281 199 282 201
rect 284 199 285 201
rect 281 205 282 207
rect 284 205 285 207
rect 301 219 302 221
rect 304 219 305 221
rect 301 225 302 227
rect 304 225 305 227
rect 221 179 222 181
rect 224 179 225 181
rect 221 185 222 187
rect 224 185 225 187
rect 241 359 242 361
rect 244 359 245 361
rect 241 365 242 367
rect 244 365 245 367
rect 441 199 442 201
rect 444 199 445 201
rect 441 205 442 207
rect 444 205 445 207
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect 161 19 162 21
rect 164 19 165 21
rect 161 25 162 27
rect 164 25 165 27
rect 161 79 162 81
rect 164 79 165 81
rect 161 85 162 87
rect 164 85 165 87
rect 161 279 162 281
rect 164 279 165 281
rect 161 285 162 287
rect 164 285 165 287
rect 41 199 42 201
rect 44 199 45 201
rect 41 205 42 207
rect 44 205 45 207
rect 201 179 202 181
rect 204 179 205 181
rect 201 185 202 187
rect 204 185 205 187
rect 181 339 182 341
rect 184 339 185 341
rect 181 345 182 347
rect 184 345 185 347
rect 81 199 82 201
rect 84 199 85 201
rect 81 205 82 207
rect 84 205 85 207
rect 301 259 302 261
rect 304 259 305 261
rect 301 265 302 267
rect 304 265 305 267
rect 201 379 202 381
rect 204 379 205 381
rect 201 385 202 387
rect 204 385 205 387
rect 221 279 222 281
rect 224 279 225 281
rect 221 285 222 287
rect 224 285 225 287
rect 261 419 262 421
rect 264 419 265 421
rect 261 425 262 427
rect 264 425 265 427
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect 61 339 62 341
rect 64 339 65 341
rect 61 345 62 347
rect 64 345 65 347
rect 121 259 122 261
rect 124 259 125 261
rect 121 265 122 267
rect 124 265 125 267
rect 141 99 142 101
rect 144 99 145 101
rect 141 105 142 107
rect 144 105 145 107
rect 341 319 342 321
rect 344 319 345 321
rect 341 325 342 327
rect 344 325 345 327
rect 141 19 142 21
rect 144 19 145 21
rect 141 25 142 27
rect 144 25 145 27
rect 61 259 62 261
rect 64 259 65 261
rect 61 265 62 267
rect 64 265 65 267
rect 241 439 242 441
rect 244 439 245 441
rect 241 445 242 447
rect 244 445 245 447
rect 241 119 242 121
rect 244 119 245 121
rect 241 125 242 127
rect 244 125 245 127
rect 141 179 142 181
rect 144 179 145 181
rect 141 185 142 187
rect 144 185 145 187
rect 281 39 282 41
rect 284 39 285 41
rect 281 45 282 47
rect 284 45 285 47
rect 361 199 362 201
rect 364 199 365 201
rect 361 205 362 207
rect 364 205 365 207
rect 341 379 342 381
rect 344 379 345 381
rect 341 385 342 387
rect 344 385 345 387
rect 1 279 2 281
rect 4 279 5 281
rect 1 285 2 287
rect 4 285 5 287
rect 301 79 302 81
rect 304 79 305 81
rect 301 85 302 87
rect 304 85 305 87
rect 281 359 282 361
rect 284 359 285 361
rect 281 365 282 367
rect 284 365 285 367
rect 121 299 122 301
rect 124 299 125 301
rect 121 305 122 307
rect 124 305 125 307
rect 221 119 222 121
rect 224 119 225 121
rect 221 125 222 127
rect 224 125 225 127
rect 161 39 162 41
rect 164 39 165 41
rect 161 45 162 47
rect 164 45 165 47
rect 261 -1 262 1
rect 264 -1 265 1
rect 261 5 262 7
rect 264 5 265 7
rect 241 179 242 181
rect 244 179 245 181
rect 241 185 242 187
rect 244 185 245 187
rect 201 339 202 341
rect 204 339 205 341
rect 201 345 202 347
rect 204 345 205 347
rect 341 159 342 161
rect 344 159 345 161
rect 341 165 342 167
rect 344 165 345 167
rect 121 39 122 41
rect 124 39 125 41
rect 121 45 122 47
rect 124 45 125 47
rect 301 239 302 241
rect 304 239 305 241
rect 301 245 302 247
rect 304 245 305 247
rect 281 419 282 421
rect 284 419 285 421
rect 281 425 282 427
rect 284 425 285 427
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect 181 239 182 241
rect 184 239 185 241
rect 181 245 182 247
rect 184 245 185 247
rect 261 59 262 61
rect 264 59 265 61
rect 261 65 262 67
rect 264 65 265 67
rect 261 279 262 281
rect 264 279 265 281
rect 261 285 262 287
rect 264 285 265 287
rect 321 119 322 121
rect 324 119 325 121
rect 321 125 322 127
rect 324 125 325 127
rect 301 199 302 201
rect 304 199 305 201
rect 301 205 302 207
rect 304 205 305 207
rect 321 339 322 341
rect 324 339 325 341
rect 321 345 322 347
rect 324 345 325 347
rect 241 139 242 141
rect 244 139 245 141
rect 241 145 242 147
rect 244 145 245 147
rect 61 139 62 141
rect 64 139 65 141
rect 61 145 62 147
rect 64 145 65 147
rect 361 119 362 121
rect 364 119 365 121
rect 361 125 362 127
rect 364 125 365 127
rect 201 239 202 241
rect 204 239 205 241
rect 201 245 202 247
rect 204 245 205 247
rect 341 179 342 181
rect 344 179 345 181
rect 341 185 342 187
rect 344 185 345 187
rect 61 179 62 181
rect 64 179 65 181
rect 61 185 62 187
rect 64 185 65 187
rect 181 39 182 41
rect 184 39 185 41
rect 181 45 182 47
rect 184 45 185 47
rect 201 459 202 461
rect 204 459 205 461
rect 201 465 202 467
rect 204 465 205 467
rect 341 99 342 101
rect 344 99 345 101
rect 341 105 342 107
rect 344 105 345 107
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect 261 79 262 81
rect 264 79 265 81
rect 261 85 262 87
rect 264 85 265 87
rect 181 59 182 61
rect 184 59 185 61
rect 181 65 182 67
rect 184 65 185 67
rect 21 139 22 141
rect 24 139 25 141
rect 21 145 22 147
rect 24 145 25 147
rect 41 119 42 121
rect 44 119 45 121
rect 41 125 42 127
rect 44 125 45 127
rect 381 259 382 261
rect 384 259 385 261
rect 381 265 382 267
rect 384 265 385 267
rect 221 419 222 421
rect 224 419 225 421
rect 221 425 222 427
rect 224 425 225 427
rect 301 119 302 121
rect 304 119 305 121
rect 301 125 302 127
rect 304 125 305 127
rect 221 39 222 41
rect 224 39 225 41
rect 221 45 222 47
rect 224 45 225 47
rect 201 159 202 161
rect 204 159 205 161
rect 201 165 202 167
rect 204 165 205 167
rect 21 119 22 121
rect 24 119 25 121
rect 21 125 22 127
rect 24 125 25 127
rect 161 239 162 241
rect 164 239 165 241
rect 161 245 162 247
rect 164 245 165 247
rect 321 419 322 421
rect 324 419 325 421
rect 321 425 322 427
rect 324 425 325 427
rect 221 19 222 21
rect 224 19 225 21
rect 221 25 222 27
rect 224 25 225 27
rect 221 79 222 81
rect 224 79 225 81
rect 221 85 222 87
rect 224 85 225 87
rect 321 159 322 161
rect 324 159 325 161
rect 321 165 322 167
rect 324 165 325 167
rect 141 199 142 201
rect 144 199 145 201
rect 141 205 142 207
rect 144 205 145 207
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect 401 219 402 221
rect 404 219 405 221
rect 401 225 402 227
rect 404 225 405 227
rect 181 279 182 281
rect 184 279 185 281
rect 181 285 182 287
rect 184 285 185 287
rect 201 299 202 301
rect 204 299 205 301
rect 201 305 202 307
rect 204 305 205 307
rect 301 439 302 441
rect 304 439 305 441
rect 301 445 302 447
rect 304 445 305 447
rect 101 259 102 261
rect 104 259 105 261
rect 101 265 102 267
rect 104 265 105 267
rect 341 79 342 81
rect 344 79 345 81
rect 341 85 342 87
rect 344 85 345 87
rect 161 -1 162 1
rect 164 -1 165 1
rect 161 5 162 7
rect 164 5 165 7
rect 41 299 42 301
rect 44 299 45 301
rect 41 305 42 307
rect 44 305 45 307
rect 141 259 142 261
rect 144 259 145 261
rect 141 265 142 267
rect 144 265 145 267
rect 241 19 242 21
rect 244 19 245 21
rect 241 25 242 27
rect 244 25 245 27
rect 141 379 142 381
rect 144 379 145 381
rect 141 385 142 387
rect 144 385 145 387
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect 241 79 242 81
rect 244 79 245 81
rect 241 85 242 87
rect 244 85 245 87
rect 41 259 42 261
rect 44 259 45 261
rect 41 265 42 267
rect 44 265 45 267
rect 121 99 122 101
rect 124 99 125 101
rect 121 105 122 107
rect 124 105 125 107
rect 321 79 322 81
rect 324 79 325 81
rect 321 85 322 87
rect 324 85 325 87
rect 321 179 322 181
rect 324 179 325 181
rect 321 185 322 187
rect 324 185 325 187
rect 281 339 282 341
rect 284 339 285 341
rect 281 345 282 347
rect 284 345 285 347
rect 221 399 222 401
rect 224 399 225 401
rect 221 405 222 407
rect 224 405 225 407
rect 101 179 102 181
rect 104 179 105 181
rect 101 185 102 187
rect 104 185 105 187
rect 181 399 182 401
rect 184 399 185 401
rect 181 405 182 407
rect 184 405 185 407
rect 181 439 182 441
rect 184 439 185 441
rect 181 445 182 447
rect 184 445 185 447
rect 221 379 222 381
rect 224 379 225 381
rect 221 385 222 387
rect 224 385 225 387
rect 401 119 402 121
rect 404 119 405 121
rect 401 125 402 127
rect 404 125 405 127
rect 381 199 382 201
rect 384 199 385 201
rect 381 205 382 207
rect 384 205 385 207
rect 261 179 262 181
rect 264 179 265 181
rect 261 185 262 187
rect 264 185 265 187
rect 341 119 342 121
rect 344 119 345 121
rect 341 125 342 127
rect 344 125 345 127
rect 161 399 162 401
rect 164 399 165 401
rect 161 405 162 407
rect 164 405 165 407
rect 1 99 2 101
rect 4 99 5 101
rect 1 105 2 107
rect 4 105 5 107
rect 81 59 82 61
rect 84 59 85 61
rect 81 65 82 67
rect 84 65 85 67
rect 1 159 2 161
rect 4 159 5 161
rect 1 165 2 167
rect 4 165 5 167
rect 281 459 282 461
rect 284 459 285 461
rect 281 465 282 467
rect 284 465 285 467
rect 161 139 162 141
rect 164 139 165 141
rect 161 145 162 147
rect 164 145 165 147
rect 181 299 182 301
rect 184 299 185 301
rect 181 305 182 307
rect 184 305 185 307
rect 421 179 422 181
rect 424 179 425 181
rect 421 185 422 187
rect 424 185 425 187
rect 141 339 142 341
rect 144 339 145 341
rect 141 345 142 347
rect 144 345 145 347
rect 361 319 362 321
rect 364 319 365 321
rect 361 325 362 327
rect 364 325 365 327
rect 281 119 282 121
rect 284 119 285 121
rect 281 125 282 127
rect 284 125 285 127
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect 141 359 142 361
rect 144 359 145 361
rect 141 365 142 367
rect 144 365 145 367
rect 181 99 182 101
rect 184 99 185 101
rect 181 105 182 107
rect 184 105 185 107
rect 101 39 102 41
rect 104 39 105 41
rect 101 45 102 47
rect 104 45 105 47
rect 101 59 102 61
rect 104 59 105 61
rect 101 65 102 67
rect 104 65 105 67
rect 261 259 262 261
rect 264 259 265 261
rect 261 265 262 267
rect 264 265 265 267
rect 241 379 242 381
rect 244 379 245 381
rect 241 385 242 387
rect 244 385 245 387
rect 21 239 22 241
rect 24 239 25 241
rect 21 245 22 247
rect 24 245 25 247
rect 61 119 62 121
rect 64 119 65 121
rect 61 125 62 127
rect 64 125 65 127
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect 181 259 182 261
rect 184 259 185 261
rect 181 265 182 267
rect 184 265 185 267
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect 221 319 222 321
rect 224 319 225 321
rect 221 325 222 327
rect 224 325 225 327
rect 161 419 162 421
rect 164 419 165 421
rect 161 425 162 427
rect 164 425 165 427
rect 321 439 322 441
rect 324 439 325 441
rect 321 445 322 447
rect 324 445 325 447
rect 101 119 102 121
rect 104 119 105 121
rect 101 125 102 127
rect 104 125 105 127
rect 281 219 282 221
rect 284 219 285 221
rect 281 225 282 227
rect 284 225 285 227
rect 141 419 142 421
rect 144 419 145 421
rect 141 425 142 427
rect 144 425 145 427
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect 261 99 262 101
rect 264 99 265 101
rect 261 105 262 107
rect 264 105 265 107
rect 241 99 242 101
rect 244 99 245 101
rect 241 105 242 107
rect 244 105 245 107
rect 81 239 82 241
rect 84 239 85 241
rect 81 245 82 247
rect 84 245 85 247
rect 341 359 342 361
rect 344 359 345 361
rect 341 365 342 367
rect 344 365 345 367
rect 241 339 242 341
rect 244 339 245 341
rect 241 345 242 347
rect 244 345 245 347
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect 241 219 242 221
rect 244 219 245 221
rect 241 225 242 227
rect 244 225 245 227
rect 301 139 302 141
rect 304 139 305 141
rect 301 145 302 147
rect 304 145 305 147
rect 241 59 242 61
rect 244 59 245 61
rect 241 65 242 67
rect 244 65 245 67
rect 21 199 22 201
rect 24 199 25 201
rect 21 205 22 207
rect 24 205 25 207
rect 141 139 142 141
rect 144 139 145 141
rect 141 145 142 147
rect 144 145 145 147
rect 261 19 262 21
rect 264 19 265 21
rect 261 25 262 27
rect 264 25 265 27
rect 361 179 362 181
rect 364 179 365 181
rect 361 185 362 187
rect 364 185 365 187
rect 301 419 302 421
rect 304 419 305 421
rect 301 425 302 427
rect 304 425 305 427
rect 201 359 202 361
rect 204 359 205 361
rect 201 365 202 367
rect 204 365 205 367
rect 101 199 102 201
rect 104 199 105 201
rect 101 205 102 207
rect 104 205 105 207
rect 161 379 162 381
rect 164 379 165 381
rect 161 385 162 387
rect 164 385 165 387
rect 261 319 262 321
rect 264 319 265 321
rect 261 325 262 327
rect 264 325 265 327
rect 381 239 382 241
rect 384 239 385 241
rect 381 245 382 247
rect 384 245 385 247
rect 41 279 42 281
rect 44 279 45 281
rect 41 285 42 287
rect 44 285 45 287
rect 301 59 302 61
rect 304 59 305 61
rect 301 65 302 67
rect 304 65 305 67
rect 101 279 102 281
rect 104 279 105 281
rect 101 285 102 287
rect 104 285 105 287
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect 81 259 82 261
rect 84 259 85 261
rect 81 265 82 267
rect 84 265 85 267
rect 381 179 382 181
rect 384 179 385 181
rect 381 185 382 187
rect 384 185 385 187
rect 381 359 382 361
rect 384 359 385 361
rect 381 365 382 367
rect 384 365 385 367
rect 141 299 142 301
rect 144 299 145 301
rect 141 305 142 307
rect 144 305 145 307
rect 341 259 342 261
rect 344 259 345 261
rect 341 265 342 267
rect 344 265 345 267
rect 101 359 102 361
rect 104 359 105 361
rect 101 365 102 367
rect 104 365 105 367
rect 141 219 142 221
rect 144 219 145 221
rect 141 225 142 227
rect 144 225 145 227
rect 241 419 242 421
rect 244 419 245 421
rect 241 425 242 427
rect 244 425 245 427
<< labels >>
rlabel pdiffusion 123 323 124 324 0 Cellno = 1
rlabel pdiffusion 363 243 364 244 0 Cellno = 2
rlabel pdiffusion 143 323 144 324 0 Cellno = 3
rlabel pdiffusion 263 363 264 364 0 Cellno = 4
rlabel pdiffusion 183 383 184 384 0 Cellno = 5
rlabel pdiffusion 323 243 324 244 0 Cellno = 6
rlabel pdiffusion 83 403 84 404 0 Cellno = 7
rlabel pdiffusion 83 303 84 304 0 Cellno = 8
rlabel pdiffusion 363 163 364 164 0 Cellno = 9
rlabel pdiffusion 323 203 324 204 0 Cellno = 10
rlabel pdiffusion 323 323 324 324 0 Cellno = 11
rlabel pdiffusion 383 163 384 164 0 Cellno = 12
rlabel pdiffusion 283 403 284 404 0 Cellno = 13
rlabel pdiffusion 3 143 4 144 0 Cellno = 14
rlabel pdiffusion 103 343 104 344 0 Cellno = 15
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 16
rlabel pdiffusion 83 283 84 284 0 Cellno = 17
rlabel pdiffusion 123 363 124 364 0 Cellno = 18
rlabel pdiffusion 83 163 84 164 0 Cellno = 19
rlabel pdiffusion 323 223 324 224 0 Cellno = 20
rlabel pdiffusion 263 443 264 444 0 Cellno = 21
rlabel pdiffusion 203 283 204 284 0 Cellno = 22
rlabel pdiffusion 363 263 364 264 0 Cellno = 23
rlabel pdiffusion 403 243 404 244 0 Cellno = 24
rlabel pdiffusion 83 123 84 124 0 Cellno = 25
rlabel pdiffusion 323 403 324 404 0 Cellno = 26
rlabel pdiffusion 263 303 264 304 0 Cellno = 27
rlabel pdiffusion 163 303 164 304 0 Cellno = 28
rlabel pdiffusion 263 43 264 44 0 Cellno = 29
rlabel pdiffusion 243 263 244 264 0 Cellno = 30
rlabel pdiffusion 183 123 184 124 0 Cellno = 31
rlabel pdiffusion 43 143 44 144 0 Cellno = 32
rlabel pdiffusion 403 263 404 264 0 Cellno = 33
rlabel pdiffusion 243 303 244 304 0 Cellno = 34
rlabel pdiffusion 163 183 164 184 0 Cellno = 35
rlabel pdiffusion 263 343 264 344 0 Cellno = 36
rlabel pdiffusion 123 243 124 244 0 Cellno = 37
rlabel pdiffusion 403 163 404 164 0 Cellno = 38
rlabel pdiffusion 43 163 44 164 0 Cellno = 39
rlabel pdiffusion 283 383 284 384 0 Cellno = 40
rlabel pdiffusion 143 403 144 404 0 Cellno = 41
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 42
rlabel pdiffusion 283 103 284 104 0 Cellno = 43
rlabel pdiffusion 103 83 104 84 0 Cellno = 44
rlabel pdiffusion 403 203 404 204 0 Cellno = 45
rlabel pdiffusion 283 303 284 304 0 Cellno = 46
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 47
rlabel pdiffusion 283 443 284 444 0 Cellno = 48
rlabel pdiffusion 163 343 164 344 0 Cellno = 49
rlabel pdiffusion 103 103 104 104 0 Cellno = 50
rlabel pdiffusion 203 223 204 224 0 Cellno = 51
rlabel pdiffusion 103 323 104 324 0 Cellno = 52
rlabel pdiffusion 163 263 164 264 0 Cellno = 53
rlabel pdiffusion 123 203 124 204 0 Cellno = 54
rlabel pdiffusion 283 63 284 64 0 Cellno = 55
rlabel pdiffusion 83 323 84 324 0 Cellno = 56
rlabel pdiffusion 363 363 364 364 0 Cellno = 57
rlabel pdiffusion 203 123 204 124 0 Cellno = 58
rlabel pdiffusion 243 283 244 284 0 Cellno = 59
rlabel pdiffusion 263 223 264 224 0 Cellno = 60
rlabel pdiffusion 223 203 224 204 0 Cellno = 61
rlabel pdiffusion 263 403 264 404 0 Cellno = 62
rlabel pdiffusion 143 243 144 244 0 Cellno = 63
rlabel pdiffusion 243 163 244 164 0 Cellno = 64
rlabel pdiffusion 103 243 104 244 0 Cellno = 65
rlabel pdiffusion 163 323 164 324 0 Cellno = 66
rlabel pdiffusion 163 163 164 164 0 Cellno = 67
rlabel pdiffusion 83 363 84 364 0 Cellno = 68
rlabel pdiffusion 43 103 44 104 0 Cellno = 69
rlabel pdiffusion 203 443 204 444 0 Cellno = 70
rlabel pdiffusion 63 203 64 204 0 Cellno = 71
rlabel pdiffusion 3 183 4 184 0 Cellno = 72
rlabel pdiffusion 183 203 184 204 0 Cellno = 73
rlabel pdiffusion 303 403 304 404 0 Cellno = 74
rlabel pdiffusion 303 163 304 164 0 Cellno = 75
rlabel pdiffusion 3 223 4 224 0 Cellno = 76
rlabel pdiffusion 383 143 384 144 0 Cellno = 77
rlabel pdiffusion 83 43 84 44 0 Cellno = 78
rlabel pdiffusion 123 343 124 344 0 Cellno = 79
rlabel pdiffusion 63 303 64 304 0 Cellno = 80
rlabel pdiffusion 243 3 244 4 0 Cellno = 81
rlabel pdiffusion 283 243 284 244 0 Cellno = 82
rlabel pdiffusion 43 323 44 324 0 Cellno = 83
rlabel pdiffusion 203 103 204 104 0 Cellno = 84
rlabel pdiffusion 303 103 304 104 0 Cellno = 85
rlabel pdiffusion 323 303 324 304 0 Cellno = 86
rlabel pdiffusion 3 123 4 124 0 Cellno = 87
rlabel pdiffusion 423 243 424 244 0 Cellno = 88
rlabel pdiffusion 303 343 304 344 0 Cellno = 89
rlabel pdiffusion 163 203 164 204 0 Cellno = 90
rlabel pdiffusion 103 143 104 144 0 Cellno = 91
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 92
rlabel pdiffusion 383 283 384 284 0 Cellno = 93
rlabel pdiffusion 23 163 24 164 0 Cellno = 94
rlabel pdiffusion 123 183 124 184 0 Cellno = 95
rlabel pdiffusion 123 123 124 124 0 Cellno = 96
rlabel pdiffusion 423 203 424 204 0 Cellno = 97
rlabel pdiffusion 223 243 224 244 0 Cellno = 98
rlabel pdiffusion 243 243 244 244 0 Cellno = 99
rlabel pdiffusion 423 223 424 224 0 Cellno = 100
rlabel pdiffusion 183 423 184 424 0 Cellno = 101
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 102
rlabel pdiffusion 343 403 344 404 0 Cellno = 103
rlabel pdiffusion 83 223 84 224 0 Cellno = 104
rlabel pdiffusion 43 243 44 244 0 Cellno = 105
rlabel pdiffusion 183 363 184 364 0 Cellno = 106
rlabel pdiffusion 343 223 344 224 0 Cellno = 107
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 108
rlabel pdiffusion 283 3 284 4 0 Cellno = 109
rlabel pdiffusion 263 163 264 164 0 Cellno = 110
rlabel pdiffusion 283 323 284 324 0 Cellno = 111
rlabel pdiffusion 123 223 124 224 0 Cellno = 112
rlabel pdiffusion 63 163 64 164 0 Cellno = 113
rlabel pdiffusion 263 123 264 124 0 Cellno = 114
rlabel pdiffusion 163 103 164 104 0 Cellno = 115
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 116
rlabel pdiffusion 363 223 364 224 0 Cellno = 117
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 118
rlabel pdiffusion 103 403 104 404 0 Cellno = 119
rlabel pdiffusion 423 123 424 124 0 Cellno = 120
rlabel pdiffusion 23 183 24 184 0 Cellno = 121
rlabel pdiffusion 203 63 204 64 0 Cellno = 122
rlabel pdiffusion 83 83 84 84 0 Cellno = 123
rlabel pdiffusion 243 403 244 404 0 Cellno = 124
rlabel pdiffusion 63 243 64 244 0 Cellno = 125
rlabel pdiffusion 143 163 144 164 0 Cellno = 126
rlabel pdiffusion 303 323 304 324 0 Cellno = 127
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 128
rlabel pdiffusion 203 23 204 24 0 Cellno = 129
rlabel pdiffusion 283 23 284 24 0 Cellno = 130
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 131
rlabel pdiffusion 183 323 184 324 0 Cellno = 132
rlabel pdiffusion 223 143 224 144 0 Cellno = 133
rlabel pdiffusion 323 63 324 64 0 Cellno = 134
rlabel pdiffusion 23 223 24 224 0 Cellno = 135
rlabel pdiffusion 283 263 284 264 0 Cellno = 136
rlabel pdiffusion 143 283 144 284 0 Cellno = 137
rlabel pdiffusion 303 283 304 284 0 Cellno = 138
rlabel pdiffusion 403 183 404 184 0 Cellno = 139
rlabel pdiffusion 143 123 144 124 0 Cellno = 140
rlabel pdiffusion 123 143 124 144 0 Cellno = 141
rlabel pdiffusion 263 203 264 204 0 Cellno = 142
rlabel pdiffusion 163 223 164 224 0 Cellno = 143
rlabel pdiffusion 263 463 264 464 0 Cellno = 144
rlabel pdiffusion 123 63 124 64 0 Cellno = 145
rlabel pdiffusion 303 363 304 364 0 Cellno = 146
rlabel pdiffusion 203 143 204 144 0 Cellno = 147
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 148
rlabel pdiffusion 103 163 104 164 0 Cellno = 149
rlabel pdiffusion 243 43 244 44 0 Cellno = 150
rlabel pdiffusion 223 303 224 304 0 Cellno = 151
rlabel pdiffusion 203 83 204 84 0 Cellno = 152
rlabel pdiffusion 203 43 204 44 0 Cellno = 153
rlabel pdiffusion 323 363 324 364 0 Cellno = 154
rlabel pdiffusion 343 283 344 284 0 Cellno = 155
rlabel pdiffusion 363 103 364 104 0 Cellno = 156
rlabel pdiffusion 83 143 84 144 0 Cellno = 157
rlabel pdiffusion 63 83 64 84 0 Cellno = 158
rlabel pdiffusion 123 283 124 284 0 Cellno = 159
rlabel pdiffusion 263 243 264 244 0 Cellno = 160
rlabel pdiffusion 323 383 324 384 0 Cellno = 161
rlabel pdiffusion 163 363 164 364 0 Cellno = 162
rlabel pdiffusion 223 103 224 104 0 Cellno = 163
rlabel pdiffusion 183 83 184 84 0 Cellno = 164
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 165
rlabel pdiffusion 243 323 244 324 0 Cellno = 166
rlabel pdiffusion 303 303 304 304 0 Cellno = 167
rlabel pdiffusion 203 323 204 324 0 Cellno = 168
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 169
rlabel pdiffusion 63 323 64 324 0 Cellno = 170
rlabel pdiffusion 223 163 224 164 0 Cellno = 171
rlabel pdiffusion 83 383 84 384 0 Cellno = 172
rlabel pdiffusion 263 383 264 384 0 Cellno = 173
rlabel pdiffusion 343 343 344 344 0 Cellno = 174
rlabel pdiffusion 283 163 284 164 0 Cellno = 175
rlabel pdiffusion 23 283 24 284 0 Cellno = 176
rlabel pdiffusion 363 283 364 284 0 Cellno = 177
rlabel pdiffusion 43 223 44 224 0 Cellno = 178
rlabel pdiffusion 143 63 144 64 0 Cellno = 179
rlabel pdiffusion 183 163 184 164 0 Cellno = 180
rlabel pdiffusion 363 383 364 384 0 Cellno = 181
rlabel pdiffusion 83 183 84 184 0 Cellno = 182
rlabel pdiffusion 223 263 224 264 0 Cellno = 183
rlabel pdiffusion 343 143 344 144 0 Cellno = 184
rlabel pdiffusion 143 43 144 44 0 Cellno = 185
rlabel pdiffusion 103 383 104 384 0 Cellno = 186
rlabel pdiffusion 343 203 344 204 0 Cellno = 187
rlabel pdiffusion 323 283 324 284 0 Cellno = 188
rlabel pdiffusion 203 263 204 264 0 Cellno = 189
rlabel pdiffusion 203 403 204 404 0 Cellno = 190
rlabel pdiffusion 83 103 84 104 0 Cellno = 191
rlabel pdiffusion 63 103 64 104 0 Cellno = 192
rlabel pdiffusion 143 83 144 84 0 Cellno = 193
rlabel pdiffusion 283 143 284 144 0 Cellno = 194
rlabel pdiffusion 303 183 304 184 0 Cellno = 195
rlabel pdiffusion 343 303 344 304 0 Cellno = 196
rlabel pdiffusion 403 303 404 304 0 Cellno = 197
rlabel pdiffusion 223 363 224 364 0 Cellno = 198
rlabel pdiffusion 183 223 184 224 0 Cellno = 199
rlabel pdiffusion 163 63 164 64 0 Cellno = 200
rlabel pdiffusion 43 183 44 184 0 Cellno = 201
rlabel pdiffusion 63 283 64 284 0 Cellno = 202
rlabel pdiffusion 183 183 184 184 0 Cellno = 203
rlabel pdiffusion 163 123 164 124 0 Cellno = 204
rlabel pdiffusion 383 323 384 324 0 Cellno = 205
rlabel pdiffusion 243 203 244 204 0 Cellno = 206
rlabel pdiffusion 83 343 84 344 0 Cellno = 207
rlabel pdiffusion 363 303 364 304 0 Cellno = 208
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 209
rlabel pdiffusion 303 383 304 384 0 Cellno = 210
rlabel pdiffusion 323 263 324 264 0 Cellno = 211
rlabel pdiffusion 343 243 344 244 0 Cellno = 212
rlabel pdiffusion 123 163 124 164 0 Cellno = 213
rlabel pdiffusion 283 183 284 184 0 Cellno = 214
rlabel pdiffusion 223 343 224 344 0 Cellno = 215
rlabel pdiffusion 103 223 104 224 0 Cellno = 216
rlabel pdiffusion 183 143 184 144 0 Cellno = 217
rlabel pdiffusion 363 343 364 344 0 Cellno = 218
rlabel pdiffusion 63 223 64 224 0 Cellno = 219
rlabel pdiffusion 283 283 284 284 0 Cellno = 220
rlabel pdiffusion 323 103 324 104 0 Cellno = 221
rlabel pdiffusion 383 223 384 224 0 Cellno = 222
rlabel pdiffusion 123 83 124 84 0 Cellno = 223
rlabel pdiffusion 323 143 324 144 0 Cellno = 224
rlabel pdiffusion 3 263 4 264 0 Cellno = 225
rlabel pdiffusion 323 43 324 44 0 Cellno = 226
rlabel pdiffusion 223 223 224 224 0 Cellno = 227
rlabel pdiffusion 103 303 104 304 0 Cellno = 228
rlabel pdiffusion 283 83 284 84 0 Cellno = 229
rlabel pdiffusion 183 23 184 24 0 Cellno = 230
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 231
rlabel pdiffusion 223 63 224 64 0 Cellno = 232
rlabel pdiffusion 203 203 204 204 0 Cellno = 233
rlabel pdiffusion 263 143 264 144 0 Cellno = 234
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 235
rlabel pdiffusion 283 203 284 204 0 Cellno = 236
rlabel pdiffusion 303 223 304 224 0 Cellno = 237
rlabel pdiffusion 223 183 224 184 0 Cellno = 238
rlabel pdiffusion 243 363 244 364 0 Cellno = 239
rlabel pdiffusion 443 203 444 204 0 Cellno = 240
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 241
rlabel pdiffusion 163 23 164 24 0 Cellno = 242
rlabel pdiffusion 163 83 164 84 0 Cellno = 243
rlabel pdiffusion 163 283 164 284 0 Cellno = 244
rlabel pdiffusion 43 203 44 204 0 Cellno = 245
rlabel pdiffusion 203 183 204 184 0 Cellno = 246
rlabel pdiffusion 183 343 184 344 0 Cellno = 247
rlabel pdiffusion 83 203 84 204 0 Cellno = 248
rlabel pdiffusion 303 263 304 264 0 Cellno = 249
rlabel pdiffusion 203 383 204 384 0 Cellno = 250
rlabel pdiffusion 223 283 224 284 0 Cellno = 251
rlabel pdiffusion 263 423 264 424 0 Cellno = 252
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 253
rlabel pdiffusion 63 343 64 344 0 Cellno = 254
rlabel pdiffusion 123 263 124 264 0 Cellno = 255
rlabel pdiffusion 143 103 144 104 0 Cellno = 256
rlabel pdiffusion 343 323 344 324 0 Cellno = 257
rlabel pdiffusion 143 23 144 24 0 Cellno = 258
rlabel pdiffusion 63 263 64 264 0 Cellno = 259
rlabel pdiffusion 243 443 244 444 0 Cellno = 260
rlabel pdiffusion 243 123 244 124 0 Cellno = 261
rlabel pdiffusion 143 183 144 184 0 Cellno = 262
rlabel pdiffusion 283 43 284 44 0 Cellno = 263
rlabel pdiffusion 363 203 364 204 0 Cellno = 264
rlabel pdiffusion 343 383 344 384 0 Cellno = 265
rlabel pdiffusion 3 283 4 284 0 Cellno = 266
rlabel pdiffusion 303 83 304 84 0 Cellno = 267
rlabel pdiffusion 283 363 284 364 0 Cellno = 268
rlabel pdiffusion 123 303 124 304 0 Cellno = 269
rlabel pdiffusion 223 123 224 124 0 Cellno = 270
rlabel pdiffusion 163 43 164 44 0 Cellno = 271
rlabel pdiffusion 263 3 264 4 0 Cellno = 272
rlabel pdiffusion 243 183 244 184 0 Cellno = 273
rlabel pdiffusion 203 343 204 344 0 Cellno = 274
rlabel pdiffusion 343 163 344 164 0 Cellno = 275
rlabel pdiffusion 123 43 124 44 0 Cellno = 276
rlabel pdiffusion 303 243 304 244 0 Cellno = 277
rlabel pdiffusion 283 423 284 424 0 Cellno = 278
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 279
rlabel pdiffusion 183 243 184 244 0 Cellno = 280
rlabel pdiffusion 263 63 264 64 0 Cellno = 281
rlabel pdiffusion 263 283 264 284 0 Cellno = 282
rlabel pdiffusion 323 123 324 124 0 Cellno = 283
rlabel pdiffusion 303 203 304 204 0 Cellno = 284
rlabel pdiffusion 323 343 324 344 0 Cellno = 285
rlabel pdiffusion 243 143 244 144 0 Cellno = 286
rlabel pdiffusion 63 143 64 144 0 Cellno = 287
rlabel pdiffusion 363 123 364 124 0 Cellno = 288
rlabel pdiffusion 203 243 204 244 0 Cellno = 289
rlabel pdiffusion 343 183 344 184 0 Cellno = 290
rlabel pdiffusion 63 183 64 184 0 Cellno = 291
rlabel pdiffusion 183 43 184 44 0 Cellno = 292
rlabel pdiffusion 203 463 204 464 0 Cellno = 293
rlabel pdiffusion 343 103 344 104 0 Cellno = 294
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 295
rlabel pdiffusion 263 83 264 84 0 Cellno = 296
rlabel pdiffusion 183 63 184 64 0 Cellno = 297
rlabel pdiffusion 23 143 24 144 0 Cellno = 298
rlabel pdiffusion 43 123 44 124 0 Cellno = 299
rlabel pdiffusion 383 263 384 264 0 Cellno = 300
rlabel pdiffusion 223 423 224 424 0 Cellno = 301
rlabel pdiffusion 303 123 304 124 0 Cellno = 302
rlabel pdiffusion 223 43 224 44 0 Cellno = 303
rlabel pdiffusion 203 163 204 164 0 Cellno = 304
rlabel pdiffusion 23 123 24 124 0 Cellno = 305
rlabel pdiffusion 163 243 164 244 0 Cellno = 306
rlabel pdiffusion 323 423 324 424 0 Cellno = 307
rlabel pdiffusion 223 23 224 24 0 Cellno = 308
rlabel pdiffusion 223 83 224 84 0 Cellno = 309
rlabel pdiffusion 323 163 324 164 0 Cellno = 310
rlabel pdiffusion 143 203 144 204 0 Cellno = 311
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 312
rlabel pdiffusion 403 223 404 224 0 Cellno = 313
rlabel pdiffusion 183 283 184 284 0 Cellno = 314
rlabel pdiffusion 203 303 204 304 0 Cellno = 315
rlabel pdiffusion 303 443 304 444 0 Cellno = 316
rlabel pdiffusion 103 263 104 264 0 Cellno = 317
rlabel pdiffusion 343 83 344 84 0 Cellno = 318
rlabel pdiffusion 163 3 164 4 0 Cellno = 319
rlabel pdiffusion 43 303 44 304 0 Cellno = 320
rlabel pdiffusion 143 263 144 264 0 Cellno = 321
rlabel pdiffusion 243 23 244 24 0 Cellno = 322
rlabel pdiffusion 143 383 144 384 0 Cellno = 323
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 324
rlabel pdiffusion 243 83 244 84 0 Cellno = 325
rlabel pdiffusion 43 263 44 264 0 Cellno = 326
rlabel pdiffusion 123 103 124 104 0 Cellno = 327
rlabel pdiffusion 323 83 324 84 0 Cellno = 328
rlabel pdiffusion 323 183 324 184 0 Cellno = 329
rlabel pdiffusion 283 343 284 344 0 Cellno = 330
rlabel pdiffusion 223 403 224 404 0 Cellno = 331
rlabel pdiffusion 103 183 104 184 0 Cellno = 332
rlabel pdiffusion 183 403 184 404 0 Cellno = 333
rlabel pdiffusion 183 443 184 444 0 Cellno = 334
rlabel pdiffusion 223 383 224 384 0 Cellno = 335
rlabel pdiffusion 403 123 404 124 0 Cellno = 336
rlabel pdiffusion 383 203 384 204 0 Cellno = 337
rlabel pdiffusion 263 183 264 184 0 Cellno = 338
rlabel pdiffusion 343 123 344 124 0 Cellno = 339
rlabel pdiffusion 163 403 164 404 0 Cellno = 340
rlabel pdiffusion 3 103 4 104 0 Cellno = 341
rlabel pdiffusion 83 63 84 64 0 Cellno = 342
rlabel pdiffusion 3 163 4 164 0 Cellno = 343
rlabel pdiffusion 283 463 284 464 0 Cellno = 344
rlabel pdiffusion 163 143 164 144 0 Cellno = 345
rlabel pdiffusion 183 303 184 304 0 Cellno = 346
rlabel pdiffusion 423 183 424 184 0 Cellno = 347
rlabel pdiffusion 143 343 144 344 0 Cellno = 348
rlabel pdiffusion 363 323 364 324 0 Cellno = 349
rlabel pdiffusion 283 123 284 124 0 Cellno = 350
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 351
rlabel pdiffusion 143 363 144 364 0 Cellno = 352
rlabel pdiffusion 183 103 184 104 0 Cellno = 353
rlabel pdiffusion 103 43 104 44 0 Cellno = 354
rlabel pdiffusion 103 63 104 64 0 Cellno = 355
rlabel pdiffusion 263 263 264 264 0 Cellno = 356
rlabel pdiffusion 243 383 244 384 0 Cellno = 357
rlabel pdiffusion 23 243 24 244 0 Cellno = 358
rlabel pdiffusion 63 123 64 124 0 Cellno = 359
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 360
rlabel pdiffusion 183 263 184 264 0 Cellno = 361
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 362
rlabel pdiffusion 223 323 224 324 0 Cellno = 363
rlabel pdiffusion 163 423 164 424 0 Cellno = 364
rlabel pdiffusion 323 443 324 444 0 Cellno = 365
rlabel pdiffusion 103 123 104 124 0 Cellno = 366
rlabel pdiffusion 283 223 284 224 0 Cellno = 367
rlabel pdiffusion 143 423 144 424 0 Cellno = 368
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 369
rlabel pdiffusion 263 103 264 104 0 Cellno = 370
rlabel pdiffusion 243 103 244 104 0 Cellno = 371
rlabel pdiffusion 83 243 84 244 0 Cellno = 372
rlabel pdiffusion 343 363 344 364 0 Cellno = 373
rlabel pdiffusion 243 343 244 344 0 Cellno = 374
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 375
rlabel pdiffusion 243 223 244 224 0 Cellno = 376
rlabel pdiffusion 303 143 304 144 0 Cellno = 377
rlabel pdiffusion 243 63 244 64 0 Cellno = 378
rlabel pdiffusion 23 203 24 204 0 Cellno = 379
rlabel pdiffusion 143 143 144 144 0 Cellno = 380
rlabel pdiffusion 263 23 264 24 0 Cellno = 381
rlabel pdiffusion 363 183 364 184 0 Cellno = 382
rlabel pdiffusion 303 423 304 424 0 Cellno = 383
rlabel pdiffusion 203 363 204 364 0 Cellno = 384
rlabel pdiffusion 103 203 104 204 0 Cellno = 385
rlabel pdiffusion 163 383 164 384 0 Cellno = 386
rlabel pdiffusion 263 323 264 324 0 Cellno = 387
rlabel pdiffusion 383 243 384 244 0 Cellno = 388
rlabel pdiffusion 43 283 44 284 0 Cellno = 389
rlabel pdiffusion 303 63 304 64 0 Cellno = 390
rlabel pdiffusion 103 283 104 284 0 Cellno = 391
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 392
rlabel pdiffusion 83 263 84 264 0 Cellno = 393
rlabel pdiffusion 383 183 384 184 0 Cellno = 394
rlabel pdiffusion 383 363 384 364 0 Cellno = 395
rlabel pdiffusion 143 303 144 304 0 Cellno = 396
rlabel pdiffusion 343 263 344 264 0 Cellno = 397
rlabel pdiffusion 103 363 104 364 0 Cellno = 398
rlabel pdiffusion 143 223 144 224 0 Cellno = 399
rlabel pdiffusion 243 423 244 424 0 Cellno = 400
<< end >>
