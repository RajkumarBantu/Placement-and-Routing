magic
tech scmos
timestamp
<< pdiffusion >>
rect 680 700 681 701
rect 682 700 683 701
rect 683 700 684 701
rect 685 700 686 701
rect 680 701 686 705
rect 680 705 681 706
rect 682 705 683 706
rect 683 705 684 706
rect 685 705 686 706
rect 580 420 581 421
rect 582 420 583 421
rect 583 420 584 421
rect 585 420 586 421
rect 580 421 586 425
rect 580 425 581 426
rect 582 425 583 426
rect 583 425 584 426
rect 585 425 586 426
rect 740 600 741 601
rect 742 600 743 601
rect 743 600 744 601
rect 745 600 746 601
rect 740 601 746 605
rect 740 605 741 606
rect 742 605 743 606
rect 743 605 744 606
rect 745 605 746 606
rect 760 520 761 521
rect 762 520 763 521
rect 763 520 764 521
rect 765 520 766 521
rect 760 521 766 525
rect 760 525 761 526
rect 762 525 763 526
rect 763 525 764 526
rect 765 525 766 526
rect 640 840 641 841
rect 642 840 643 841
rect 643 840 644 841
rect 645 840 646 841
rect 640 841 646 845
rect 640 845 641 846
rect 642 845 643 846
rect 643 845 644 846
rect 645 845 646 846
rect 640 740 641 741
rect 642 740 643 741
rect 643 740 644 741
rect 645 740 646 741
rect 640 741 646 745
rect 640 745 641 746
rect 642 745 643 746
rect 643 745 644 746
rect 645 745 646 746
rect 600 920 601 921
rect 602 920 603 921
rect 603 920 604 921
rect 605 920 606 921
rect 600 921 606 925
rect 600 925 601 926
rect 602 925 603 926
rect 603 925 604 926
rect 605 925 606 926
rect 500 800 501 801
rect 502 800 503 801
rect 503 800 504 801
rect 505 800 506 801
rect 500 801 506 805
rect 500 805 501 806
rect 502 805 503 806
rect 503 805 504 806
rect 505 805 506 806
rect 800 660 801 661
rect 802 660 803 661
rect 803 660 804 661
rect 805 660 806 661
rect 800 661 806 665
rect 800 665 801 666
rect 802 665 803 666
rect 803 665 804 666
rect 805 665 806 666
rect 480 640 481 641
rect 482 640 483 641
rect 483 640 484 641
rect 485 640 486 641
rect 480 641 486 645
rect 480 645 481 646
rect 482 645 483 646
rect 483 645 484 646
rect 485 645 486 646
rect 840 620 841 621
rect 842 620 843 621
rect 843 620 844 621
rect 845 620 846 621
rect 840 621 846 625
rect 840 625 841 626
rect 842 625 843 626
rect 843 625 844 626
rect 845 625 846 626
rect 760 660 761 661
rect 762 660 763 661
rect 763 660 764 661
rect 765 660 766 661
rect 760 661 766 665
rect 760 665 761 666
rect 762 665 763 666
rect 763 665 764 666
rect 765 665 766 666
rect 700 700 701 701
rect 702 700 703 701
rect 703 700 704 701
rect 705 700 706 701
rect 700 701 706 705
rect 700 705 701 706
rect 702 705 703 706
rect 703 705 704 706
rect 705 705 706 706
rect 520 540 521 541
rect 522 540 523 541
rect 523 540 524 541
rect 525 540 526 541
rect 520 541 526 545
rect 520 545 521 546
rect 522 545 523 546
rect 523 545 524 546
rect 525 545 526 546
rect 420 860 421 861
rect 422 860 423 861
rect 423 860 424 861
rect 425 860 426 861
rect 420 861 426 865
rect 420 865 421 866
rect 422 865 423 866
rect 423 865 424 866
rect 425 865 426 866
rect 600 900 601 901
rect 602 900 603 901
rect 603 900 604 901
rect 605 900 606 901
rect 600 901 606 905
rect 600 905 601 906
rect 602 905 603 906
rect 603 905 604 906
rect 605 905 606 906
rect 440 840 441 841
rect 442 840 443 841
rect 443 840 444 841
rect 445 840 446 841
rect 440 841 446 845
rect 440 845 441 846
rect 442 845 443 846
rect 443 845 444 846
rect 445 845 446 846
rect 680 740 681 741
rect 682 740 683 741
rect 683 740 684 741
rect 685 740 686 741
rect 680 741 686 745
rect 680 745 681 746
rect 682 745 683 746
rect 683 745 684 746
rect 685 745 686 746
rect 540 540 541 541
rect 542 540 543 541
rect 543 540 544 541
rect 545 540 546 541
rect 540 541 546 545
rect 540 545 541 546
rect 542 545 543 546
rect 543 545 544 546
rect 545 545 546 546
rect 860 740 861 741
rect 862 740 863 741
rect 863 740 864 741
rect 865 740 866 741
rect 860 741 866 745
rect 860 745 861 746
rect 862 745 863 746
rect 863 745 864 746
rect 865 745 866 746
rect 560 880 561 881
rect 562 880 563 881
rect 563 880 564 881
rect 565 880 566 881
rect 560 881 566 885
rect 560 885 561 886
rect 562 885 563 886
rect 563 885 564 886
rect 565 885 566 886
rect 560 600 561 601
rect 562 600 563 601
rect 563 600 564 601
rect 565 600 566 601
rect 560 601 566 605
rect 560 605 561 606
rect 562 605 563 606
rect 563 605 564 606
rect 565 605 566 606
rect 640 540 641 541
rect 642 540 643 541
rect 643 540 644 541
rect 645 540 646 541
rect 640 541 646 545
rect 640 545 641 546
rect 642 545 643 546
rect 643 545 644 546
rect 645 545 646 546
rect 640 800 641 801
rect 642 800 643 801
rect 643 800 644 801
rect 645 800 646 801
rect 640 801 646 805
rect 640 805 641 806
rect 642 805 643 806
rect 643 805 644 806
rect 645 805 646 806
rect 540 800 541 801
rect 542 800 543 801
rect 543 800 544 801
rect 545 800 546 801
rect 540 801 546 805
rect 540 805 541 806
rect 542 805 543 806
rect 543 805 544 806
rect 545 805 546 806
rect 580 900 581 901
rect 582 900 583 901
rect 583 900 584 901
rect 585 900 586 901
rect 580 901 586 905
rect 580 905 581 906
rect 582 905 583 906
rect 583 905 584 906
rect 585 905 586 906
rect 920 720 921 721
rect 922 720 923 721
rect 923 720 924 721
rect 925 720 926 721
rect 920 721 926 725
rect 920 725 921 726
rect 922 725 923 726
rect 923 725 924 726
rect 925 725 926 726
rect 480 760 481 761
rect 482 760 483 761
rect 483 760 484 761
rect 485 760 486 761
rect 480 761 486 765
rect 480 765 481 766
rect 482 765 483 766
rect 483 765 484 766
rect 485 765 486 766
rect 680 660 681 661
rect 682 660 683 661
rect 683 660 684 661
rect 685 660 686 661
rect 680 661 686 665
rect 680 665 681 666
rect 682 665 683 666
rect 683 665 684 666
rect 685 665 686 666
rect 680 840 681 841
rect 682 840 683 841
rect 683 840 684 841
rect 685 840 686 841
rect 680 841 686 845
rect 680 845 681 846
rect 682 845 683 846
rect 683 845 684 846
rect 685 845 686 846
rect 760 480 761 481
rect 762 480 763 481
rect 763 480 764 481
rect 765 480 766 481
rect 760 481 766 485
rect 760 485 761 486
rect 762 485 763 486
rect 763 485 764 486
rect 765 485 766 486
rect 400 840 401 841
rect 402 840 403 841
rect 403 840 404 841
rect 405 840 406 841
rect 400 841 406 845
rect 400 845 401 846
rect 402 845 403 846
rect 403 845 404 846
rect 405 845 406 846
rect 460 560 461 561
rect 462 560 463 561
rect 463 560 464 561
rect 465 560 466 561
rect 460 561 466 565
rect 460 565 461 566
rect 462 565 463 566
rect 463 565 464 566
rect 465 565 466 566
rect 440 720 441 721
rect 442 720 443 721
rect 443 720 444 721
rect 445 720 446 721
rect 440 721 446 725
rect 440 725 441 726
rect 442 725 443 726
rect 443 725 444 726
rect 445 725 446 726
rect 600 580 601 581
rect 602 580 603 581
rect 603 580 604 581
rect 605 580 606 581
rect 600 581 606 585
rect 600 585 601 586
rect 602 585 603 586
rect 603 585 604 586
rect 605 585 606 586
rect 920 700 921 701
rect 922 700 923 701
rect 923 700 924 701
rect 925 700 926 701
rect 920 701 926 705
rect 920 705 921 706
rect 922 705 923 706
rect 923 705 924 706
rect 925 705 926 706
rect 760 620 761 621
rect 762 620 763 621
rect 763 620 764 621
rect 765 620 766 621
rect 760 621 766 625
rect 760 625 761 626
rect 762 625 763 626
rect 763 625 764 626
rect 765 625 766 626
rect 700 780 701 781
rect 702 780 703 781
rect 703 780 704 781
rect 705 780 706 781
rect 700 781 706 785
rect 700 785 701 786
rect 702 785 703 786
rect 703 785 704 786
rect 705 785 706 786
rect 640 640 641 641
rect 642 640 643 641
rect 643 640 644 641
rect 645 640 646 641
rect 640 641 646 645
rect 640 645 641 646
rect 642 645 643 646
rect 643 645 644 646
rect 645 645 646 646
rect 440 700 441 701
rect 442 700 443 701
rect 443 700 444 701
rect 445 700 446 701
rect 440 701 446 705
rect 440 705 441 706
rect 442 705 443 706
rect 443 705 444 706
rect 445 705 446 706
rect 600 640 601 641
rect 602 640 603 641
rect 603 640 604 641
rect 605 640 606 641
rect 600 641 606 645
rect 600 645 601 646
rect 602 645 603 646
rect 603 645 604 646
rect 605 645 606 646
rect 720 600 721 601
rect 722 600 723 601
rect 723 600 724 601
rect 725 600 726 601
rect 720 601 726 605
rect 720 605 721 606
rect 722 605 723 606
rect 723 605 724 606
rect 725 605 726 606
rect 440 900 441 901
rect 442 900 443 901
rect 443 900 444 901
rect 445 900 446 901
rect 440 901 446 905
rect 440 905 441 906
rect 442 905 443 906
rect 443 905 444 906
rect 445 905 446 906
rect 600 520 601 521
rect 602 520 603 521
rect 603 520 604 521
rect 605 520 606 521
rect 600 521 606 525
rect 600 525 601 526
rect 602 525 603 526
rect 603 525 604 526
rect 605 525 606 526
rect 580 680 581 681
rect 582 680 583 681
rect 583 680 584 681
rect 585 680 586 681
rect 580 681 586 685
rect 580 685 581 686
rect 582 685 583 686
rect 583 685 584 686
rect 585 685 586 686
rect 720 680 721 681
rect 722 680 723 681
rect 723 680 724 681
rect 725 680 726 681
rect 720 681 726 685
rect 720 685 721 686
rect 722 685 723 686
rect 723 685 724 686
rect 725 685 726 686
rect 800 700 801 701
rect 802 700 803 701
rect 803 700 804 701
rect 805 700 806 701
rect 800 701 806 705
rect 800 705 801 706
rect 802 705 803 706
rect 803 705 804 706
rect 805 705 806 706
rect 780 580 781 581
rect 782 580 783 581
rect 783 580 784 581
rect 785 580 786 581
rect 780 581 786 585
rect 780 585 781 586
rect 782 585 783 586
rect 783 585 784 586
rect 785 585 786 586
rect 860 600 861 601
rect 862 600 863 601
rect 863 600 864 601
rect 865 600 866 601
rect 860 601 866 605
rect 860 605 861 606
rect 862 605 863 606
rect 863 605 864 606
rect 865 605 866 606
rect 500 940 501 941
rect 502 940 503 941
rect 503 940 504 941
rect 505 940 506 941
rect 500 941 506 945
rect 500 945 501 946
rect 502 945 503 946
rect 503 945 504 946
rect 505 945 506 946
rect 740 720 741 721
rect 742 720 743 721
rect 743 720 744 721
rect 745 720 746 721
rect 740 721 746 725
rect 740 725 741 726
rect 742 725 743 726
rect 743 725 744 726
rect 745 725 746 726
rect 520 760 521 761
rect 522 760 523 761
rect 523 760 524 761
rect 525 760 526 761
rect 520 761 526 765
rect 520 765 521 766
rect 522 765 523 766
rect 523 765 524 766
rect 525 765 526 766
rect 840 740 841 741
rect 842 740 843 741
rect 843 740 844 741
rect 845 740 846 741
rect 840 741 846 745
rect 840 745 841 746
rect 842 745 843 746
rect 843 745 844 746
rect 845 745 846 746
rect 700 580 701 581
rect 702 580 703 581
rect 703 580 704 581
rect 705 580 706 581
rect 700 581 706 585
rect 700 585 701 586
rect 702 585 703 586
rect 703 585 704 586
rect 705 585 706 586
rect 580 540 581 541
rect 582 540 583 541
rect 583 540 584 541
rect 585 540 586 541
rect 580 541 586 545
rect 580 545 581 546
rect 582 545 583 546
rect 583 545 584 546
rect 585 545 586 546
rect 780 760 781 761
rect 782 760 783 761
rect 783 760 784 761
rect 785 760 786 761
rect 780 761 786 765
rect 780 765 781 766
rect 782 765 783 766
rect 783 765 784 766
rect 785 765 786 766
rect 600 840 601 841
rect 602 840 603 841
rect 603 840 604 841
rect 605 840 606 841
rect 600 841 606 845
rect 600 845 601 846
rect 602 845 603 846
rect 603 845 604 846
rect 605 845 606 846
rect 660 440 661 441
rect 662 440 663 441
rect 663 440 664 441
rect 665 440 666 441
rect 660 441 666 445
rect 660 445 661 446
rect 662 445 663 446
rect 663 445 664 446
rect 665 445 666 446
rect 780 640 781 641
rect 782 640 783 641
rect 783 640 784 641
rect 785 640 786 641
rect 780 641 786 645
rect 780 645 781 646
rect 782 645 783 646
rect 783 645 784 646
rect 785 645 786 646
rect 520 680 521 681
rect 522 680 523 681
rect 523 680 524 681
rect 525 680 526 681
rect 520 681 526 685
rect 520 685 521 686
rect 522 685 523 686
rect 523 685 524 686
rect 525 685 526 686
rect 340 680 341 681
rect 342 680 343 681
rect 343 680 344 681
rect 345 680 346 681
rect 340 681 346 685
rect 340 685 341 686
rect 342 685 343 686
rect 343 685 344 686
rect 345 685 346 686
rect 480 660 481 661
rect 482 660 483 661
rect 483 660 484 661
rect 485 660 486 661
rect 480 661 486 665
rect 480 665 481 666
rect 482 665 483 666
rect 483 665 484 666
rect 485 665 486 666
rect 600 980 601 981
rect 602 980 603 981
rect 603 980 604 981
rect 605 980 606 981
rect 600 981 606 985
rect 600 985 601 986
rect 602 985 603 986
rect 603 985 604 986
rect 605 985 606 986
rect 680 600 681 601
rect 682 600 683 601
rect 683 600 684 601
rect 685 600 686 601
rect 680 601 686 605
rect 680 605 681 606
rect 682 605 683 606
rect 683 605 684 606
rect 685 605 686 606
rect 680 900 681 901
rect 682 900 683 901
rect 683 900 684 901
rect 685 900 686 901
rect 680 901 686 905
rect 680 905 681 906
rect 682 905 683 906
rect 683 905 684 906
rect 685 905 686 906
rect 820 900 821 901
rect 822 900 823 901
rect 823 900 824 901
rect 825 900 826 901
rect 820 901 826 905
rect 820 905 821 906
rect 822 905 823 906
rect 823 905 824 906
rect 825 905 826 906
rect 660 780 661 781
rect 662 780 663 781
rect 663 780 664 781
rect 665 780 666 781
rect 660 781 666 785
rect 660 785 661 786
rect 662 785 663 786
rect 663 785 664 786
rect 665 785 666 786
rect 680 860 681 861
rect 682 860 683 861
rect 683 860 684 861
rect 685 860 686 861
rect 680 861 686 865
rect 680 865 681 866
rect 682 865 683 866
rect 683 865 684 866
rect 685 865 686 866
rect 660 880 661 881
rect 662 880 663 881
rect 663 880 664 881
rect 665 880 666 881
rect 660 881 666 885
rect 660 885 661 886
rect 662 885 663 886
rect 663 885 664 886
rect 665 885 666 886
rect 340 700 341 701
rect 342 700 343 701
rect 343 700 344 701
rect 345 700 346 701
rect 340 701 346 705
rect 340 705 341 706
rect 342 705 343 706
rect 343 705 344 706
rect 345 705 346 706
rect 540 560 541 561
rect 542 560 543 561
rect 543 560 544 561
rect 545 560 546 561
rect 540 561 546 565
rect 540 565 541 566
rect 542 565 543 566
rect 543 565 544 566
rect 545 565 546 566
rect 380 860 381 861
rect 382 860 383 861
rect 383 860 384 861
rect 385 860 386 861
rect 380 861 386 865
rect 380 865 381 866
rect 382 865 383 866
rect 383 865 384 866
rect 385 865 386 866
rect 720 740 721 741
rect 722 740 723 741
rect 723 740 724 741
rect 725 740 726 741
rect 720 741 726 745
rect 720 745 721 746
rect 722 745 723 746
rect 723 745 724 746
rect 725 745 726 746
rect 520 740 521 741
rect 522 740 523 741
rect 523 740 524 741
rect 525 740 526 741
rect 520 741 526 745
rect 520 745 521 746
rect 522 745 523 746
rect 523 745 524 746
rect 525 745 526 746
rect 620 880 621 881
rect 622 880 623 881
rect 623 880 624 881
rect 625 880 626 881
rect 620 881 626 885
rect 620 885 621 886
rect 622 885 623 886
rect 623 885 624 886
rect 625 885 626 886
rect 620 380 621 381
rect 622 380 623 381
rect 623 380 624 381
rect 625 380 626 381
rect 620 381 626 385
rect 620 385 621 386
rect 622 385 623 386
rect 623 385 624 386
rect 625 385 626 386
rect 660 620 661 621
rect 662 620 663 621
rect 663 620 664 621
rect 665 620 666 621
rect 660 621 666 625
rect 660 625 661 626
rect 662 625 663 626
rect 663 625 664 626
rect 665 625 666 626
rect 760 700 761 701
rect 762 700 763 701
rect 763 700 764 701
rect 765 700 766 701
rect 760 701 766 705
rect 760 705 761 706
rect 762 705 763 706
rect 763 705 764 706
rect 765 705 766 706
rect 860 500 861 501
rect 862 500 863 501
rect 863 500 864 501
rect 865 500 866 501
rect 860 501 866 505
rect 860 505 861 506
rect 862 505 863 506
rect 863 505 864 506
rect 865 505 866 506
rect 500 840 501 841
rect 502 840 503 841
rect 503 840 504 841
rect 505 840 506 841
rect 500 841 506 845
rect 500 845 501 846
rect 502 845 503 846
rect 503 845 504 846
rect 505 845 506 846
rect 700 480 701 481
rect 702 480 703 481
rect 703 480 704 481
rect 705 480 706 481
rect 700 481 706 485
rect 700 485 701 486
rect 702 485 703 486
rect 703 485 704 486
rect 705 485 706 486
rect 520 560 521 561
rect 522 560 523 561
rect 523 560 524 561
rect 525 560 526 561
rect 520 561 526 565
rect 520 565 521 566
rect 522 565 523 566
rect 523 565 524 566
rect 525 565 526 566
rect 960 680 961 681
rect 962 680 963 681
rect 963 680 964 681
rect 965 680 966 681
rect 960 681 966 685
rect 960 685 961 686
rect 962 685 963 686
rect 963 685 964 686
rect 965 685 966 686
rect 440 560 441 561
rect 442 560 443 561
rect 443 560 444 561
rect 445 560 446 561
rect 440 561 446 565
rect 440 565 441 566
rect 442 565 443 566
rect 443 565 444 566
rect 445 565 446 566
rect 480 780 481 781
rect 482 780 483 781
rect 483 780 484 781
rect 485 780 486 781
rect 480 781 486 785
rect 480 785 481 786
rect 482 785 483 786
rect 483 785 484 786
rect 485 785 486 786
rect 480 880 481 881
rect 482 880 483 881
rect 483 880 484 881
rect 485 880 486 881
rect 480 881 486 885
rect 480 885 481 886
rect 482 885 483 886
rect 483 885 484 886
rect 485 885 486 886
rect 660 680 661 681
rect 662 680 663 681
rect 663 680 664 681
rect 665 680 666 681
rect 660 681 666 685
rect 660 685 661 686
rect 662 685 663 686
rect 663 685 664 686
rect 665 685 666 686
rect 640 460 641 461
rect 642 460 643 461
rect 643 460 644 461
rect 645 460 646 461
rect 640 461 646 465
rect 640 465 641 466
rect 642 465 643 466
rect 643 465 644 466
rect 645 465 646 466
rect 840 840 841 841
rect 842 840 843 841
rect 843 840 844 841
rect 845 840 846 841
rect 840 841 846 845
rect 840 845 841 846
rect 842 845 843 846
rect 843 845 844 846
rect 845 845 846 846
rect 620 680 621 681
rect 622 680 623 681
rect 623 680 624 681
rect 625 680 626 681
rect 620 681 626 685
rect 620 685 621 686
rect 622 685 623 686
rect 623 685 624 686
rect 625 685 626 686
rect 920 780 921 781
rect 922 780 923 781
rect 923 780 924 781
rect 925 780 926 781
rect 920 781 926 785
rect 920 785 921 786
rect 922 785 923 786
rect 923 785 924 786
rect 925 785 926 786
rect 440 640 441 641
rect 442 640 443 641
rect 443 640 444 641
rect 445 640 446 641
rect 440 641 446 645
rect 440 645 441 646
rect 442 645 443 646
rect 443 645 444 646
rect 445 645 446 646
rect 920 800 921 801
rect 922 800 923 801
rect 923 800 924 801
rect 925 800 926 801
rect 920 801 926 805
rect 920 805 921 806
rect 922 805 923 806
rect 923 805 924 806
rect 925 805 926 806
rect 380 600 381 601
rect 382 600 383 601
rect 383 600 384 601
rect 385 600 386 601
rect 380 601 386 605
rect 380 605 381 606
rect 382 605 383 606
rect 383 605 384 606
rect 385 605 386 606
rect 800 820 801 821
rect 802 820 803 821
rect 803 820 804 821
rect 805 820 806 821
rect 800 821 806 825
rect 800 825 801 826
rect 802 825 803 826
rect 803 825 804 826
rect 805 825 806 826
rect 460 920 461 921
rect 462 920 463 921
rect 463 920 464 921
rect 465 920 466 921
rect 460 921 466 925
rect 460 925 461 926
rect 462 925 463 926
rect 463 925 464 926
rect 465 925 466 926
rect 360 540 361 541
rect 362 540 363 541
rect 363 540 364 541
rect 365 540 366 541
rect 360 541 366 545
rect 360 545 361 546
rect 362 545 363 546
rect 363 545 364 546
rect 365 545 366 546
rect 660 560 661 561
rect 662 560 663 561
rect 663 560 664 561
rect 665 560 666 561
rect 660 561 666 565
rect 660 565 661 566
rect 662 565 663 566
rect 663 565 664 566
rect 665 565 666 566
rect 640 480 641 481
rect 642 480 643 481
rect 643 480 644 481
rect 645 480 646 481
rect 640 481 646 485
rect 640 485 641 486
rect 642 485 643 486
rect 643 485 644 486
rect 645 485 646 486
rect 740 620 741 621
rect 742 620 743 621
rect 743 620 744 621
rect 745 620 746 621
rect 740 621 746 625
rect 740 625 741 626
rect 742 625 743 626
rect 743 625 744 626
rect 745 625 746 626
rect 660 900 661 901
rect 662 900 663 901
rect 663 900 664 901
rect 665 900 666 901
rect 660 901 666 905
rect 660 905 661 906
rect 662 905 663 906
rect 663 905 664 906
rect 665 905 666 906
rect 800 480 801 481
rect 802 480 803 481
rect 803 480 804 481
rect 805 480 806 481
rect 800 481 806 485
rect 800 485 801 486
rect 802 485 803 486
rect 803 485 804 486
rect 805 485 806 486
rect 800 720 801 721
rect 802 720 803 721
rect 803 720 804 721
rect 805 720 806 721
rect 800 721 806 725
rect 800 725 801 726
rect 802 725 803 726
rect 803 725 804 726
rect 805 725 806 726
rect 460 620 461 621
rect 462 620 463 621
rect 463 620 464 621
rect 465 620 466 621
rect 460 621 466 625
rect 460 625 461 626
rect 462 625 463 626
rect 463 625 464 626
rect 465 625 466 626
rect 560 540 561 541
rect 562 540 563 541
rect 563 540 564 541
rect 565 540 566 541
rect 560 541 566 545
rect 560 545 561 546
rect 562 545 563 546
rect 563 545 564 546
rect 565 545 566 546
rect 620 720 621 721
rect 622 720 623 721
rect 623 720 624 721
rect 625 720 626 721
rect 620 721 626 725
rect 620 725 621 726
rect 622 725 623 726
rect 623 725 624 726
rect 625 725 626 726
rect 800 800 801 801
rect 802 800 803 801
rect 803 800 804 801
rect 805 800 806 801
rect 800 801 806 805
rect 800 805 801 806
rect 802 805 803 806
rect 803 805 804 806
rect 805 805 806 806
rect 600 600 601 601
rect 602 600 603 601
rect 603 600 604 601
rect 605 600 606 601
rect 600 601 606 605
rect 600 605 601 606
rect 602 605 603 606
rect 603 605 604 606
rect 605 605 606 606
rect 920 840 921 841
rect 922 840 923 841
rect 923 840 924 841
rect 925 840 926 841
rect 920 841 926 845
rect 920 845 921 846
rect 922 845 923 846
rect 923 845 924 846
rect 925 845 926 846
rect 480 540 481 541
rect 482 540 483 541
rect 483 540 484 541
rect 485 540 486 541
rect 480 541 486 545
rect 480 545 481 546
rect 482 545 483 546
rect 483 545 484 546
rect 485 545 486 546
rect 920 560 921 561
rect 922 560 923 561
rect 923 560 924 561
rect 925 560 926 561
rect 920 561 926 565
rect 920 565 921 566
rect 922 565 923 566
rect 923 565 924 566
rect 925 565 926 566
rect 640 700 641 701
rect 642 700 643 701
rect 643 700 644 701
rect 645 700 646 701
rect 640 701 646 705
rect 640 705 641 706
rect 642 705 643 706
rect 643 705 644 706
rect 645 705 646 706
rect 640 520 641 521
rect 642 520 643 521
rect 643 520 644 521
rect 645 520 646 521
rect 640 521 646 525
rect 640 525 641 526
rect 642 525 643 526
rect 643 525 644 526
rect 645 525 646 526
rect 920 680 921 681
rect 922 680 923 681
rect 923 680 924 681
rect 925 680 926 681
rect 920 681 926 685
rect 920 685 921 686
rect 922 685 923 686
rect 923 685 924 686
rect 925 685 926 686
rect 620 760 621 761
rect 622 760 623 761
rect 623 760 624 761
rect 625 760 626 761
rect 620 761 626 765
rect 620 765 621 766
rect 622 765 623 766
rect 623 765 624 766
rect 625 765 626 766
rect 420 740 421 741
rect 422 740 423 741
rect 423 740 424 741
rect 425 740 426 741
rect 420 741 426 745
rect 420 745 421 746
rect 422 745 423 746
rect 423 745 424 746
rect 425 745 426 746
rect 800 520 801 521
rect 802 520 803 521
rect 803 520 804 521
rect 805 520 806 521
rect 800 521 806 525
rect 800 525 801 526
rect 802 525 803 526
rect 803 525 804 526
rect 805 525 806 526
rect 720 460 721 461
rect 722 460 723 461
rect 723 460 724 461
rect 725 460 726 461
rect 720 461 726 465
rect 720 465 721 466
rect 722 465 723 466
rect 723 465 724 466
rect 725 465 726 466
rect 920 580 921 581
rect 922 580 923 581
rect 923 580 924 581
rect 925 580 926 581
rect 920 581 926 585
rect 920 585 921 586
rect 922 585 923 586
rect 923 585 924 586
rect 925 585 926 586
rect 560 780 561 781
rect 562 780 563 781
rect 563 780 564 781
rect 565 780 566 781
rect 560 781 566 785
rect 560 785 561 786
rect 562 785 563 786
rect 563 785 564 786
rect 565 785 566 786
rect 500 380 501 381
rect 502 380 503 381
rect 503 380 504 381
rect 505 380 506 381
rect 500 381 506 385
rect 500 385 501 386
rect 502 385 503 386
rect 503 385 504 386
rect 505 385 506 386
rect 940 600 941 601
rect 942 600 943 601
rect 943 600 944 601
rect 945 600 946 601
rect 940 601 946 605
rect 940 605 941 606
rect 942 605 943 606
rect 943 605 944 606
rect 945 605 946 606
rect 420 540 421 541
rect 422 540 423 541
rect 423 540 424 541
rect 425 540 426 541
rect 420 541 426 545
rect 420 545 421 546
rect 422 545 423 546
rect 423 545 424 546
rect 425 545 426 546
rect 940 620 941 621
rect 942 620 943 621
rect 943 620 944 621
rect 945 620 946 621
rect 940 621 946 625
rect 940 625 941 626
rect 942 625 943 626
rect 943 625 944 626
rect 945 625 946 626
rect 560 720 561 721
rect 562 720 563 721
rect 563 720 564 721
rect 565 720 566 721
rect 560 721 566 725
rect 560 725 561 726
rect 562 725 563 726
rect 563 725 564 726
rect 565 725 566 726
rect 460 860 461 861
rect 462 860 463 861
rect 463 860 464 861
rect 465 860 466 861
rect 460 861 466 865
rect 460 865 461 866
rect 462 865 463 866
rect 463 865 464 866
rect 465 865 466 866
rect 560 820 561 821
rect 562 820 563 821
rect 563 820 564 821
rect 565 820 566 821
rect 560 821 566 825
rect 560 825 561 826
rect 562 825 563 826
rect 563 825 564 826
rect 565 825 566 826
rect 740 640 741 641
rect 742 640 743 641
rect 743 640 744 641
rect 745 640 746 641
rect 740 641 746 645
rect 740 645 741 646
rect 742 645 743 646
rect 743 645 744 646
rect 745 645 746 646
rect 760 880 761 881
rect 762 880 763 881
rect 763 880 764 881
rect 765 880 766 881
rect 760 881 766 885
rect 760 885 761 886
rect 762 885 763 886
rect 763 885 764 886
rect 765 885 766 886
rect 480 680 481 681
rect 482 680 483 681
rect 483 680 484 681
rect 485 680 486 681
rect 480 681 486 685
rect 480 685 481 686
rect 482 685 483 686
rect 483 685 484 686
rect 485 685 486 686
rect 840 940 841 941
rect 842 940 843 941
rect 843 940 844 941
rect 845 940 846 941
rect 840 941 846 945
rect 840 945 841 946
rect 842 945 843 946
rect 843 945 844 946
rect 845 945 846 946
rect 860 460 861 461
rect 862 460 863 461
rect 863 460 864 461
rect 865 460 866 461
rect 860 461 866 465
rect 860 465 861 466
rect 862 465 863 466
rect 863 465 864 466
rect 865 465 866 466
rect 660 600 661 601
rect 662 600 663 601
rect 663 600 664 601
rect 665 600 666 601
rect 660 601 666 605
rect 660 605 661 606
rect 662 605 663 606
rect 663 605 664 606
rect 665 605 666 606
rect 480 480 481 481
rect 482 480 483 481
rect 483 480 484 481
rect 485 480 486 481
rect 480 481 486 485
rect 480 485 481 486
rect 482 485 483 486
rect 483 485 484 486
rect 485 485 486 486
rect 720 520 721 521
rect 722 520 723 521
rect 723 520 724 521
rect 725 520 726 521
rect 720 521 726 525
rect 720 525 721 526
rect 722 525 723 526
rect 723 525 724 526
rect 725 525 726 526
rect 500 580 501 581
rect 502 580 503 581
rect 503 580 504 581
rect 505 580 506 581
rect 500 581 506 585
rect 500 585 501 586
rect 502 585 503 586
rect 503 585 504 586
rect 505 585 506 586
rect 360 840 361 841
rect 362 840 363 841
rect 363 840 364 841
rect 365 840 366 841
rect 360 841 366 845
rect 360 845 361 846
rect 362 845 363 846
rect 363 845 364 846
rect 365 845 366 846
rect 360 820 361 821
rect 362 820 363 821
rect 363 820 364 821
rect 365 820 366 821
rect 360 821 366 825
rect 360 825 361 826
rect 362 825 363 826
rect 363 825 364 826
rect 365 825 366 826
rect 740 520 741 521
rect 742 520 743 521
rect 743 520 744 521
rect 745 520 746 521
rect 740 521 746 525
rect 740 525 741 526
rect 742 525 743 526
rect 743 525 744 526
rect 745 525 746 526
rect 840 780 841 781
rect 842 780 843 781
rect 843 780 844 781
rect 845 780 846 781
rect 840 781 846 785
rect 840 785 841 786
rect 842 785 843 786
rect 843 785 844 786
rect 845 785 846 786
rect 380 620 381 621
rect 382 620 383 621
rect 383 620 384 621
rect 385 620 386 621
rect 380 621 386 625
rect 380 625 381 626
rect 382 625 383 626
rect 383 625 384 626
rect 385 625 386 626
rect 480 840 481 841
rect 482 840 483 841
rect 483 840 484 841
rect 485 840 486 841
rect 480 841 486 845
rect 480 845 481 846
rect 482 845 483 846
rect 483 845 484 846
rect 485 845 486 846
rect 560 480 561 481
rect 562 480 563 481
rect 563 480 564 481
rect 565 480 566 481
rect 560 481 566 485
rect 560 485 561 486
rect 562 485 563 486
rect 563 485 564 486
rect 565 485 566 486
rect 440 680 441 681
rect 442 680 443 681
rect 443 680 444 681
rect 445 680 446 681
rect 440 681 446 685
rect 440 685 441 686
rect 442 685 443 686
rect 443 685 444 686
rect 445 685 446 686
rect 500 700 501 701
rect 502 700 503 701
rect 503 700 504 701
rect 505 700 506 701
rect 500 701 506 705
rect 500 705 501 706
rect 502 705 503 706
rect 503 705 504 706
rect 505 705 506 706
rect 520 840 521 841
rect 522 840 523 841
rect 523 840 524 841
rect 525 840 526 841
rect 520 841 526 845
rect 520 845 521 846
rect 522 845 523 846
rect 523 845 524 846
rect 525 845 526 846
rect 540 640 541 641
rect 542 640 543 641
rect 543 640 544 641
rect 545 640 546 641
rect 540 641 546 645
rect 540 645 541 646
rect 542 645 543 646
rect 543 645 544 646
rect 545 645 546 646
rect 800 560 801 561
rect 802 560 803 561
rect 803 560 804 561
rect 805 560 806 561
rect 800 561 806 565
rect 800 565 801 566
rect 802 565 803 566
rect 803 565 804 566
rect 805 565 806 566
rect 560 520 561 521
rect 562 520 563 521
rect 563 520 564 521
rect 565 520 566 521
rect 560 521 566 525
rect 560 525 561 526
rect 562 525 563 526
rect 563 525 564 526
rect 565 525 566 526
rect 580 700 581 701
rect 582 700 583 701
rect 583 700 584 701
rect 585 700 586 701
rect 580 701 586 705
rect 580 705 581 706
rect 582 705 583 706
rect 583 705 584 706
rect 585 705 586 706
rect 600 800 601 801
rect 602 800 603 801
rect 603 800 604 801
rect 605 800 606 801
rect 600 801 606 805
rect 600 805 601 806
rect 602 805 603 806
rect 603 805 604 806
rect 605 805 606 806
rect 820 880 821 881
rect 822 880 823 881
rect 823 880 824 881
rect 825 880 826 881
rect 820 881 826 885
rect 820 885 821 886
rect 822 885 823 886
rect 823 885 824 886
rect 825 885 826 886
rect 760 780 761 781
rect 762 780 763 781
rect 763 780 764 781
rect 765 780 766 781
rect 760 781 766 785
rect 760 785 761 786
rect 762 785 763 786
rect 763 785 764 786
rect 765 785 766 786
rect 620 960 621 961
rect 622 960 623 961
rect 623 960 624 961
rect 625 960 626 961
rect 620 961 626 965
rect 620 965 621 966
rect 622 965 623 966
rect 623 965 624 966
rect 625 965 626 966
rect 480 700 481 701
rect 482 700 483 701
rect 483 700 484 701
rect 485 700 486 701
rect 480 701 486 705
rect 480 705 481 706
rect 482 705 483 706
rect 483 705 484 706
rect 485 705 486 706
rect 500 440 501 441
rect 502 440 503 441
rect 503 440 504 441
rect 505 440 506 441
rect 500 441 506 445
rect 500 445 501 446
rect 502 445 503 446
rect 503 445 504 446
rect 505 445 506 446
rect 520 640 521 641
rect 522 640 523 641
rect 523 640 524 641
rect 525 640 526 641
rect 520 641 526 645
rect 520 645 521 646
rect 522 645 523 646
rect 523 645 524 646
rect 525 645 526 646
rect 760 680 761 681
rect 762 680 763 681
rect 763 680 764 681
rect 765 680 766 681
rect 760 681 766 685
rect 760 685 761 686
rect 762 685 763 686
rect 763 685 764 686
rect 765 685 766 686
rect 540 820 541 821
rect 542 820 543 821
rect 543 820 544 821
rect 545 820 546 821
rect 540 821 546 825
rect 540 825 541 826
rect 542 825 543 826
rect 543 825 544 826
rect 545 825 546 826
rect 560 380 561 381
rect 562 380 563 381
rect 563 380 564 381
rect 565 380 566 381
rect 560 381 566 385
rect 560 385 561 386
rect 562 385 563 386
rect 563 385 564 386
rect 565 385 566 386
rect 860 780 861 781
rect 862 780 863 781
rect 863 780 864 781
rect 865 780 866 781
rect 860 781 866 785
rect 860 785 861 786
rect 862 785 863 786
rect 863 785 864 786
rect 865 785 866 786
rect 660 460 661 461
rect 662 460 663 461
rect 663 460 664 461
rect 665 460 666 461
rect 660 461 666 465
rect 660 465 661 466
rect 662 465 663 466
rect 663 465 664 466
rect 665 465 666 466
rect 680 300 681 301
rect 682 300 683 301
rect 683 300 684 301
rect 685 300 686 301
rect 680 301 686 305
rect 680 305 681 306
rect 682 305 683 306
rect 683 305 684 306
rect 685 305 686 306
rect 640 620 641 621
rect 642 620 643 621
rect 643 620 644 621
rect 645 620 646 621
rect 640 621 646 625
rect 640 625 641 626
rect 642 625 643 626
rect 643 625 644 626
rect 645 625 646 626
rect 560 660 561 661
rect 562 660 563 661
rect 563 660 564 661
rect 565 660 566 661
rect 560 661 566 665
rect 560 665 561 666
rect 562 665 563 666
rect 563 665 564 666
rect 565 665 566 666
rect 360 600 361 601
rect 362 600 363 601
rect 363 600 364 601
rect 365 600 366 601
rect 360 601 366 605
rect 360 605 361 606
rect 362 605 363 606
rect 363 605 364 606
rect 365 605 366 606
rect 640 1020 641 1021
rect 642 1020 643 1021
rect 643 1020 644 1021
rect 645 1020 646 1021
rect 640 1021 646 1025
rect 640 1025 641 1026
rect 642 1025 643 1026
rect 643 1025 644 1026
rect 645 1025 646 1026
rect 720 820 721 821
rect 722 820 723 821
rect 723 820 724 821
rect 725 820 726 821
rect 720 821 726 825
rect 720 825 721 826
rect 722 825 723 826
rect 723 825 724 826
rect 725 825 726 826
rect 760 720 761 721
rect 762 720 763 721
rect 763 720 764 721
rect 765 720 766 721
rect 760 721 766 725
rect 760 725 761 726
rect 762 725 763 726
rect 763 725 764 726
rect 765 725 766 726
rect 660 800 661 801
rect 662 800 663 801
rect 663 800 664 801
rect 665 800 666 801
rect 660 801 666 805
rect 660 805 661 806
rect 662 805 663 806
rect 663 805 664 806
rect 665 805 666 806
rect 560 680 561 681
rect 562 680 563 681
rect 563 680 564 681
rect 565 680 566 681
rect 560 681 566 685
rect 560 685 561 686
rect 562 685 563 686
rect 563 685 564 686
rect 565 685 566 686
rect 460 740 461 741
rect 462 740 463 741
rect 463 740 464 741
rect 465 740 466 741
rect 460 741 466 745
rect 460 745 461 746
rect 462 745 463 746
rect 463 745 464 746
rect 465 745 466 746
rect 740 320 741 321
rect 742 320 743 321
rect 743 320 744 321
rect 745 320 746 321
rect 740 321 746 325
rect 740 325 741 326
rect 742 325 743 326
rect 743 325 744 326
rect 745 325 746 326
rect 700 520 701 521
rect 702 520 703 521
rect 703 520 704 521
rect 705 520 706 521
rect 700 521 706 525
rect 700 525 701 526
rect 702 525 703 526
rect 703 525 704 526
rect 705 525 706 526
rect 500 720 501 721
rect 502 720 503 721
rect 503 720 504 721
rect 505 720 506 721
rect 500 721 506 725
rect 500 725 501 726
rect 502 725 503 726
rect 503 725 504 726
rect 505 725 506 726
rect 700 900 701 901
rect 702 900 703 901
rect 703 900 704 901
rect 705 900 706 901
rect 700 901 706 905
rect 700 905 701 906
rect 702 905 703 906
rect 703 905 704 906
rect 705 905 706 906
rect 960 580 961 581
rect 962 580 963 581
rect 963 580 964 581
rect 965 580 966 581
rect 960 581 966 585
rect 960 585 961 586
rect 962 585 963 586
rect 963 585 964 586
rect 965 585 966 586
rect 740 960 741 961
rect 742 960 743 961
rect 743 960 744 961
rect 745 960 746 961
rect 740 961 746 965
rect 740 965 741 966
rect 742 965 743 966
rect 743 965 744 966
rect 745 965 746 966
rect 600 1040 601 1041
rect 602 1040 603 1041
rect 603 1040 604 1041
rect 605 1040 606 1041
rect 600 1041 606 1045
rect 600 1045 601 1046
rect 602 1045 603 1046
rect 603 1045 604 1046
rect 605 1045 606 1046
rect 760 940 761 941
rect 762 940 763 941
rect 763 940 764 941
rect 765 940 766 941
rect 760 941 766 945
rect 760 945 761 946
rect 762 945 763 946
rect 763 945 764 946
rect 765 945 766 946
rect 800 640 801 641
rect 802 640 803 641
rect 803 640 804 641
rect 805 640 806 641
rect 800 641 806 645
rect 800 645 801 646
rect 802 645 803 646
rect 803 645 804 646
rect 805 645 806 646
rect 320 760 321 761
rect 322 760 323 761
rect 323 760 324 761
rect 325 760 326 761
rect 320 761 326 765
rect 320 765 321 766
rect 322 765 323 766
rect 323 765 324 766
rect 325 765 326 766
rect 820 600 821 601
rect 822 600 823 601
rect 823 600 824 601
rect 825 600 826 601
rect 820 601 826 605
rect 820 605 821 606
rect 822 605 823 606
rect 823 605 824 606
rect 825 605 826 606
rect 720 300 721 301
rect 722 300 723 301
rect 723 300 724 301
rect 725 300 726 301
rect 720 301 726 305
rect 720 305 721 306
rect 722 305 723 306
rect 723 305 724 306
rect 725 305 726 306
rect 680 460 681 461
rect 682 460 683 461
rect 683 460 684 461
rect 685 460 686 461
rect 680 461 686 465
rect 680 465 681 466
rect 682 465 683 466
rect 683 465 684 466
rect 685 465 686 466
rect 820 560 821 561
rect 822 560 823 561
rect 823 560 824 561
rect 825 560 826 561
rect 820 561 826 565
rect 820 565 821 566
rect 822 565 823 566
rect 823 565 824 566
rect 825 565 826 566
rect 720 800 721 801
rect 722 800 723 801
rect 723 800 724 801
rect 725 800 726 801
rect 720 801 726 805
rect 720 805 721 806
rect 722 805 723 806
rect 723 805 724 806
rect 725 805 726 806
rect 620 920 621 921
rect 622 920 623 921
rect 623 920 624 921
rect 625 920 626 921
rect 620 921 626 925
rect 620 925 621 926
rect 622 925 623 926
rect 623 925 624 926
rect 625 925 626 926
rect 360 800 361 801
rect 362 800 363 801
rect 363 800 364 801
rect 365 800 366 801
rect 360 801 366 805
rect 360 805 361 806
rect 362 805 363 806
rect 363 805 364 806
rect 365 805 366 806
rect 540 760 541 761
rect 542 760 543 761
rect 543 760 544 761
rect 545 760 546 761
rect 540 761 546 765
rect 540 765 541 766
rect 542 765 543 766
rect 543 765 544 766
rect 545 765 546 766
rect 480 500 481 501
rect 482 500 483 501
rect 483 500 484 501
rect 485 500 486 501
rect 480 501 486 505
rect 480 505 481 506
rect 482 505 483 506
rect 483 505 484 506
rect 485 505 486 506
rect 620 560 621 561
rect 622 560 623 561
rect 623 560 624 561
rect 625 560 626 561
rect 620 561 626 565
rect 620 565 621 566
rect 622 565 623 566
rect 623 565 624 566
rect 625 565 626 566
rect 700 1020 701 1021
rect 702 1020 703 1021
rect 703 1020 704 1021
rect 705 1020 706 1021
rect 700 1021 706 1025
rect 700 1025 701 1026
rect 702 1025 703 1026
rect 703 1025 704 1026
rect 705 1025 706 1026
rect 860 920 861 921
rect 862 920 863 921
rect 863 920 864 921
rect 865 920 866 921
rect 860 921 866 925
rect 860 925 861 926
rect 862 925 863 926
rect 863 925 864 926
rect 865 925 866 926
rect 860 760 861 761
rect 862 760 863 761
rect 863 760 864 761
rect 865 760 866 761
rect 860 761 866 765
rect 860 765 861 766
rect 862 765 863 766
rect 863 765 864 766
rect 865 765 866 766
rect 980 680 981 681
rect 982 680 983 681
rect 983 680 984 681
rect 985 680 986 681
rect 980 681 986 685
rect 980 685 981 686
rect 982 685 983 686
rect 983 685 984 686
rect 985 685 986 686
rect 420 840 421 841
rect 422 840 423 841
rect 423 840 424 841
rect 425 840 426 841
rect 420 841 426 845
rect 420 845 421 846
rect 422 845 423 846
rect 423 845 424 846
rect 425 845 426 846
rect 780 840 781 841
rect 782 840 783 841
rect 783 840 784 841
rect 785 840 786 841
rect 780 841 786 845
rect 780 845 781 846
rect 782 845 783 846
rect 783 845 784 846
rect 785 845 786 846
rect 840 460 841 461
rect 842 460 843 461
rect 843 460 844 461
rect 845 460 846 461
rect 840 461 846 465
rect 840 465 841 466
rect 842 465 843 466
rect 843 465 844 466
rect 845 465 846 466
rect 500 780 501 781
rect 502 780 503 781
rect 503 780 504 781
rect 505 780 506 781
rect 500 781 506 785
rect 500 785 501 786
rect 502 785 503 786
rect 503 785 504 786
rect 505 785 506 786
rect 580 600 581 601
rect 582 600 583 601
rect 583 600 584 601
rect 585 600 586 601
rect 580 601 586 605
rect 580 605 581 606
rect 582 605 583 606
rect 583 605 584 606
rect 585 605 586 606
rect 700 320 701 321
rect 702 320 703 321
rect 703 320 704 321
rect 705 320 706 321
rect 700 321 706 325
rect 700 325 701 326
rect 702 325 703 326
rect 703 325 704 326
rect 705 325 706 326
rect 560 360 561 361
rect 562 360 563 361
rect 563 360 564 361
rect 565 360 566 361
rect 560 361 566 365
rect 560 365 561 366
rect 562 365 563 366
rect 563 365 564 366
rect 565 365 566 366
rect 780 900 781 901
rect 782 900 783 901
rect 783 900 784 901
rect 785 900 786 901
rect 780 901 786 905
rect 780 905 781 906
rect 782 905 783 906
rect 783 905 784 906
rect 785 905 786 906
rect 480 440 481 441
rect 482 440 483 441
rect 483 440 484 441
rect 485 440 486 441
rect 480 441 486 445
rect 480 445 481 446
rect 482 445 483 446
rect 483 445 484 446
rect 485 445 486 446
rect 800 540 801 541
rect 802 540 803 541
rect 803 540 804 541
rect 805 540 806 541
rect 800 541 806 545
rect 800 545 801 546
rect 802 545 803 546
rect 803 545 804 546
rect 805 545 806 546
rect 760 360 761 361
rect 762 360 763 361
rect 763 360 764 361
rect 765 360 766 361
rect 760 361 766 365
rect 760 365 761 366
rect 762 365 763 366
rect 763 365 764 366
rect 765 365 766 366
rect 620 480 621 481
rect 622 480 623 481
rect 623 480 624 481
rect 625 480 626 481
rect 620 481 626 485
rect 620 485 621 486
rect 622 485 623 486
rect 623 485 624 486
rect 625 485 626 486
rect 840 680 841 681
rect 842 680 843 681
rect 843 680 844 681
rect 845 680 846 681
rect 840 681 846 685
rect 840 685 841 686
rect 842 685 843 686
rect 843 685 844 686
rect 845 685 846 686
rect 560 740 561 741
rect 562 740 563 741
rect 563 740 564 741
rect 565 740 566 741
rect 560 741 566 745
rect 560 745 561 746
rect 562 745 563 746
rect 563 745 564 746
rect 565 745 566 746
rect 900 620 901 621
rect 902 620 903 621
rect 903 620 904 621
rect 905 620 906 621
rect 900 621 906 625
rect 900 625 901 626
rect 902 625 903 626
rect 903 625 904 626
rect 905 625 906 626
rect 440 480 441 481
rect 442 480 443 481
rect 443 480 444 481
rect 445 480 446 481
rect 440 481 446 485
rect 440 485 441 486
rect 442 485 443 486
rect 443 485 444 486
rect 445 485 446 486
rect 760 400 761 401
rect 762 400 763 401
rect 763 400 764 401
rect 765 400 766 401
rect 760 401 766 405
rect 760 405 761 406
rect 762 405 763 406
rect 763 405 764 406
rect 765 405 766 406
rect 540 720 541 721
rect 542 720 543 721
rect 543 720 544 721
rect 545 720 546 721
rect 540 721 546 725
rect 540 725 541 726
rect 542 725 543 726
rect 543 725 544 726
rect 545 725 546 726
rect 660 820 661 821
rect 662 820 663 821
rect 663 820 664 821
rect 665 820 666 821
rect 660 821 666 825
rect 660 825 661 826
rect 662 825 663 826
rect 663 825 664 826
rect 665 825 666 826
rect 400 640 401 641
rect 402 640 403 641
rect 403 640 404 641
rect 405 640 406 641
rect 400 641 406 645
rect 400 645 401 646
rect 402 645 403 646
rect 403 645 404 646
rect 405 645 406 646
rect 740 1020 741 1021
rect 742 1020 743 1021
rect 743 1020 744 1021
rect 745 1020 746 1021
rect 740 1021 746 1025
rect 740 1025 741 1026
rect 742 1025 743 1026
rect 743 1025 744 1026
rect 745 1025 746 1026
rect 540 1000 541 1001
rect 542 1000 543 1001
rect 543 1000 544 1001
rect 545 1000 546 1001
rect 540 1001 546 1005
rect 540 1005 541 1006
rect 542 1005 543 1006
rect 543 1005 544 1006
rect 545 1005 546 1006
rect 780 400 781 401
rect 782 400 783 401
rect 783 400 784 401
rect 785 400 786 401
rect 780 401 786 405
rect 780 405 781 406
rect 782 405 783 406
rect 783 405 784 406
rect 785 405 786 406
rect 660 1040 661 1041
rect 662 1040 663 1041
rect 663 1040 664 1041
rect 665 1040 666 1041
rect 660 1041 666 1045
rect 660 1045 661 1046
rect 662 1045 663 1046
rect 663 1045 664 1046
rect 665 1045 666 1046
rect 600 1060 601 1061
rect 602 1060 603 1061
rect 603 1060 604 1061
rect 605 1060 606 1061
rect 600 1061 606 1065
rect 600 1065 601 1066
rect 602 1065 603 1066
rect 603 1065 604 1066
rect 605 1065 606 1066
rect 480 740 481 741
rect 482 740 483 741
rect 483 740 484 741
rect 485 740 486 741
rect 480 741 486 745
rect 480 745 481 746
rect 482 745 483 746
rect 483 745 484 746
rect 485 745 486 746
rect 460 640 461 641
rect 462 640 463 641
rect 463 640 464 641
rect 465 640 466 641
rect 460 641 466 645
rect 460 645 461 646
rect 462 645 463 646
rect 463 645 464 646
rect 465 645 466 646
rect 460 900 461 901
rect 462 900 463 901
rect 463 900 464 901
rect 465 900 466 901
rect 460 901 466 905
rect 460 905 461 906
rect 462 905 463 906
rect 463 905 464 906
rect 465 905 466 906
rect 580 460 581 461
rect 582 460 583 461
rect 583 460 584 461
rect 585 460 586 461
rect 580 461 586 465
rect 580 465 581 466
rect 582 465 583 466
rect 583 465 584 466
rect 585 465 586 466
rect 640 400 641 401
rect 642 400 643 401
rect 643 400 644 401
rect 645 400 646 401
rect 640 401 646 405
rect 640 405 641 406
rect 642 405 643 406
rect 643 405 644 406
rect 645 405 646 406
rect 960 760 961 761
rect 962 760 963 761
rect 963 760 964 761
rect 965 760 966 761
rect 960 761 966 765
rect 960 765 961 766
rect 962 765 963 766
rect 963 765 964 766
rect 965 765 966 766
rect 560 960 561 961
rect 562 960 563 961
rect 563 960 564 961
rect 565 960 566 961
rect 560 961 566 965
rect 560 965 561 966
rect 562 965 563 966
rect 563 965 564 966
rect 565 965 566 966
rect 680 260 681 261
rect 682 260 683 261
rect 683 260 684 261
rect 685 260 686 261
rect 680 261 686 265
rect 680 265 681 266
rect 682 265 683 266
rect 683 265 684 266
rect 685 265 686 266
rect 560 580 561 581
rect 562 580 563 581
rect 563 580 564 581
rect 565 580 566 581
rect 560 581 566 585
rect 560 585 561 586
rect 562 585 563 586
rect 563 585 564 586
rect 565 585 566 586
rect 680 920 681 921
rect 682 920 683 921
rect 683 920 684 921
rect 685 920 686 921
rect 680 921 686 925
rect 680 925 681 926
rect 682 925 683 926
rect 683 925 684 926
rect 685 925 686 926
rect 500 960 501 961
rect 502 960 503 961
rect 503 960 504 961
rect 505 960 506 961
rect 500 961 506 965
rect 500 965 501 966
rect 502 965 503 966
rect 503 965 504 966
rect 505 965 506 966
rect 620 320 621 321
rect 622 320 623 321
rect 623 320 624 321
rect 625 320 626 321
rect 620 321 626 325
rect 620 325 621 326
rect 622 325 623 326
rect 623 325 624 326
rect 625 325 626 326
rect 600 380 601 381
rect 602 380 603 381
rect 603 380 604 381
rect 605 380 606 381
rect 600 381 606 385
rect 600 385 601 386
rect 602 385 603 386
rect 603 385 604 386
rect 605 385 606 386
rect 880 480 881 481
rect 882 480 883 481
rect 883 480 884 481
rect 885 480 886 481
rect 880 481 886 485
rect 880 485 881 486
rect 882 485 883 486
rect 883 485 884 486
rect 885 485 886 486
rect 1000 780 1001 781
rect 1002 780 1003 781
rect 1003 780 1004 781
rect 1005 780 1006 781
rect 1000 781 1006 785
rect 1000 785 1001 786
rect 1002 785 1003 786
rect 1003 785 1004 786
rect 1005 785 1006 786
rect 260 720 261 721
rect 262 720 263 721
rect 263 720 264 721
rect 265 720 266 721
rect 260 721 266 725
rect 260 725 261 726
rect 262 725 263 726
rect 263 725 264 726
rect 265 725 266 726
rect 560 420 561 421
rect 562 420 563 421
rect 563 420 564 421
rect 565 420 566 421
rect 560 421 566 425
rect 560 425 561 426
rect 562 425 563 426
rect 563 425 564 426
rect 565 425 566 426
rect 260 740 261 741
rect 262 740 263 741
rect 263 740 264 741
rect 265 740 266 741
rect 260 741 266 745
rect 260 745 261 746
rect 262 745 263 746
rect 263 745 264 746
rect 265 745 266 746
rect 860 840 861 841
rect 862 840 863 841
rect 863 840 864 841
rect 865 840 866 841
rect 860 841 866 845
rect 860 845 861 846
rect 862 845 863 846
rect 863 845 864 846
rect 865 845 866 846
rect 460 720 461 721
rect 462 720 463 721
rect 463 720 464 721
rect 465 720 466 721
rect 460 721 466 725
rect 460 725 461 726
rect 462 725 463 726
rect 463 725 464 726
rect 465 725 466 726
rect 640 720 641 721
rect 642 720 643 721
rect 643 720 644 721
rect 645 720 646 721
rect 640 721 646 725
rect 640 725 641 726
rect 642 725 643 726
rect 643 725 644 726
rect 645 725 646 726
rect 720 360 721 361
rect 722 360 723 361
rect 723 360 724 361
rect 725 360 726 361
rect 720 361 726 365
rect 720 365 721 366
rect 722 365 723 366
rect 723 365 724 366
rect 725 365 726 366
rect 800 460 801 461
rect 802 460 803 461
rect 803 460 804 461
rect 805 460 806 461
rect 800 461 806 465
rect 800 465 801 466
rect 802 465 803 466
rect 803 465 804 466
rect 805 465 806 466
rect 780 880 781 881
rect 782 880 783 881
rect 783 880 784 881
rect 785 880 786 881
rect 780 881 786 885
rect 780 885 781 886
rect 782 885 783 886
rect 783 885 784 886
rect 785 885 786 886
rect 900 880 901 881
rect 902 880 903 881
rect 903 880 904 881
rect 905 880 906 881
rect 900 881 906 885
rect 900 885 901 886
rect 902 885 903 886
rect 903 885 904 886
rect 905 885 906 886
rect 780 460 781 461
rect 782 460 783 461
rect 783 460 784 461
rect 785 460 786 461
rect 780 461 786 465
rect 780 465 781 466
rect 782 465 783 466
rect 783 465 784 466
rect 785 465 786 466
rect 620 1040 621 1041
rect 622 1040 623 1041
rect 623 1040 624 1041
rect 625 1040 626 1041
rect 620 1041 626 1045
rect 620 1045 621 1046
rect 622 1045 623 1046
rect 623 1045 624 1046
rect 625 1045 626 1046
rect 680 680 681 681
rect 682 680 683 681
rect 683 680 684 681
rect 685 680 686 681
rect 680 681 686 685
rect 680 685 681 686
rect 682 685 683 686
rect 683 685 684 686
rect 685 685 686 686
rect 780 540 781 541
rect 782 540 783 541
rect 783 540 784 541
rect 785 540 786 541
rect 780 541 786 545
rect 780 545 781 546
rect 782 545 783 546
rect 783 545 784 546
rect 785 545 786 546
rect 700 960 701 961
rect 702 960 703 961
rect 703 960 704 961
rect 705 960 706 961
rect 700 961 706 965
rect 700 965 701 966
rect 702 965 703 966
rect 703 965 704 966
rect 705 965 706 966
rect 620 980 621 981
rect 622 980 623 981
rect 623 980 624 981
rect 625 980 626 981
rect 620 981 626 985
rect 620 985 621 986
rect 622 985 623 986
rect 623 985 624 986
rect 625 985 626 986
rect 720 640 721 641
rect 722 640 723 641
rect 723 640 724 641
rect 725 640 726 641
rect 720 641 726 645
rect 720 645 721 646
rect 722 645 723 646
rect 723 645 724 646
rect 725 645 726 646
rect 700 740 701 741
rect 702 740 703 741
rect 703 740 704 741
rect 705 740 706 741
rect 700 741 706 745
rect 700 745 701 746
rect 702 745 703 746
rect 703 745 704 746
rect 705 745 706 746
rect 580 1020 581 1021
rect 582 1020 583 1021
rect 583 1020 584 1021
rect 585 1020 586 1021
rect 580 1021 586 1025
rect 580 1025 581 1026
rect 582 1025 583 1026
rect 583 1025 584 1026
rect 585 1025 586 1026
rect 260 640 261 641
rect 262 640 263 641
rect 263 640 264 641
rect 265 640 266 641
rect 260 641 266 645
rect 260 645 261 646
rect 262 645 263 646
rect 263 645 264 646
rect 265 645 266 646
rect 500 920 501 921
rect 502 920 503 921
rect 503 920 504 921
rect 505 920 506 921
rect 500 921 506 925
rect 500 925 501 926
rect 502 925 503 926
rect 503 925 504 926
rect 505 925 506 926
rect 740 460 741 461
rect 742 460 743 461
rect 743 460 744 461
rect 745 460 746 461
rect 740 461 746 465
rect 740 465 741 466
rect 742 465 743 466
rect 743 465 744 466
rect 745 465 746 466
rect 280 740 281 741
rect 282 740 283 741
rect 283 740 284 741
rect 285 740 286 741
rect 280 741 286 745
rect 280 745 281 746
rect 282 745 283 746
rect 283 745 284 746
rect 285 745 286 746
rect 340 800 341 801
rect 342 800 343 801
rect 343 800 344 801
rect 345 800 346 801
rect 340 801 346 805
rect 340 805 341 806
rect 342 805 343 806
rect 343 805 344 806
rect 345 805 346 806
rect 620 400 621 401
rect 622 400 623 401
rect 623 400 624 401
rect 625 400 626 401
rect 620 401 626 405
rect 620 405 621 406
rect 622 405 623 406
rect 623 405 624 406
rect 625 405 626 406
rect 780 440 781 441
rect 782 440 783 441
rect 783 440 784 441
rect 785 440 786 441
rect 780 441 786 445
rect 780 445 781 446
rect 782 445 783 446
rect 783 445 784 446
rect 785 445 786 446
rect 360 640 361 641
rect 362 640 363 641
rect 363 640 364 641
rect 365 640 366 641
rect 360 641 366 645
rect 360 645 361 646
rect 362 645 363 646
rect 363 645 364 646
rect 365 645 366 646
rect 400 660 401 661
rect 402 660 403 661
rect 403 660 404 661
rect 405 660 406 661
rect 400 661 406 665
rect 400 665 401 666
rect 402 665 403 666
rect 403 665 404 666
rect 405 665 406 666
rect 520 920 521 921
rect 522 920 523 921
rect 523 920 524 921
rect 525 920 526 921
rect 520 921 526 925
rect 520 925 521 926
rect 522 925 523 926
rect 523 925 524 926
rect 525 925 526 926
rect 720 660 721 661
rect 722 660 723 661
rect 723 660 724 661
rect 725 660 726 661
rect 720 661 726 665
rect 720 665 721 666
rect 722 665 723 666
rect 723 665 724 666
rect 725 665 726 666
rect 980 760 981 761
rect 982 760 983 761
rect 983 760 984 761
rect 985 760 986 761
rect 980 761 986 765
rect 980 765 981 766
rect 982 765 983 766
rect 983 765 984 766
rect 985 765 986 766
rect 900 840 901 841
rect 902 840 903 841
rect 903 840 904 841
rect 905 840 906 841
rect 900 841 906 845
rect 900 845 901 846
rect 902 845 903 846
rect 903 845 904 846
rect 905 845 906 846
rect 600 340 601 341
rect 602 340 603 341
rect 603 340 604 341
rect 605 340 606 341
rect 600 341 606 345
rect 600 345 601 346
rect 602 345 603 346
rect 603 345 604 346
rect 605 345 606 346
rect 980 560 981 561
rect 982 560 983 561
rect 983 560 984 561
rect 985 560 986 561
rect 980 561 986 565
rect 980 565 981 566
rect 982 565 983 566
rect 983 565 984 566
rect 985 565 986 566
rect 680 640 681 641
rect 682 640 683 641
rect 683 640 684 641
rect 685 640 686 641
rect 680 641 686 645
rect 680 645 681 646
rect 682 645 683 646
rect 683 645 684 646
rect 685 645 686 646
rect 360 580 361 581
rect 362 580 363 581
rect 363 580 364 581
rect 365 580 366 581
rect 360 581 366 585
rect 360 585 361 586
rect 362 585 363 586
rect 363 585 364 586
rect 365 585 366 586
rect 600 680 601 681
rect 602 680 603 681
rect 603 680 604 681
rect 605 680 606 681
rect 600 681 606 685
rect 600 685 601 686
rect 602 685 603 686
rect 603 685 604 686
rect 605 685 606 686
rect 920 860 921 861
rect 922 860 923 861
rect 923 860 924 861
rect 925 860 926 861
rect 920 861 926 865
rect 920 865 921 866
rect 922 865 923 866
rect 923 865 924 866
rect 925 865 926 866
rect 320 700 321 701
rect 322 700 323 701
rect 323 700 324 701
rect 325 700 326 701
rect 320 701 326 705
rect 320 705 321 706
rect 322 705 323 706
rect 323 705 324 706
rect 325 705 326 706
rect 580 780 581 781
rect 582 780 583 781
rect 583 780 584 781
rect 585 780 586 781
rect 580 781 586 785
rect 580 785 581 786
rect 582 785 583 786
rect 583 785 584 786
rect 585 785 586 786
rect 700 680 701 681
rect 702 680 703 681
rect 703 680 704 681
rect 705 680 706 681
rect 700 681 706 685
rect 700 685 701 686
rect 702 685 703 686
rect 703 685 704 686
rect 705 685 706 686
rect 720 960 721 961
rect 722 960 723 961
rect 723 960 724 961
rect 725 960 726 961
rect 720 961 726 965
rect 720 965 721 966
rect 722 965 723 966
rect 723 965 724 966
rect 725 965 726 966
rect 340 740 341 741
rect 342 740 343 741
rect 343 740 344 741
rect 345 740 346 741
rect 340 741 346 745
rect 340 745 341 746
rect 342 745 343 746
rect 343 745 344 746
rect 345 745 346 746
rect 600 480 601 481
rect 602 480 603 481
rect 603 480 604 481
rect 605 480 606 481
rect 600 481 606 485
rect 600 485 601 486
rect 602 485 603 486
rect 603 485 604 486
rect 605 485 606 486
rect 560 340 561 341
rect 562 340 563 341
rect 563 340 564 341
rect 565 340 566 341
rect 560 341 566 345
rect 560 345 561 346
rect 562 345 563 346
rect 563 345 564 346
rect 565 345 566 346
rect 700 800 701 801
rect 702 800 703 801
rect 703 800 704 801
rect 705 800 706 801
rect 700 801 706 805
rect 700 805 701 806
rect 702 805 703 806
rect 703 805 704 806
rect 705 805 706 806
rect 940 580 941 581
rect 942 580 943 581
rect 943 580 944 581
rect 945 580 946 581
rect 940 581 946 585
rect 940 585 941 586
rect 942 585 943 586
rect 943 585 944 586
rect 945 585 946 586
rect 480 460 481 461
rect 482 460 483 461
rect 483 460 484 461
rect 485 460 486 461
rect 480 461 486 465
rect 480 465 481 466
rect 482 465 483 466
rect 483 465 484 466
rect 485 465 486 466
rect 420 480 421 481
rect 422 480 423 481
rect 423 480 424 481
rect 425 480 426 481
rect 420 481 426 485
rect 420 485 421 486
rect 422 485 423 486
rect 423 485 424 486
rect 425 485 426 486
rect 480 520 481 521
rect 482 520 483 521
rect 483 520 484 521
rect 485 520 486 521
rect 480 521 486 525
rect 480 525 481 526
rect 482 525 483 526
rect 483 525 484 526
rect 485 525 486 526
rect 640 280 641 281
rect 642 280 643 281
rect 643 280 644 281
rect 645 280 646 281
rect 640 281 646 285
rect 640 285 641 286
rect 642 285 643 286
rect 643 285 644 286
rect 645 285 646 286
rect 880 600 881 601
rect 882 600 883 601
rect 883 600 884 601
rect 885 600 886 601
rect 880 601 886 605
rect 880 605 881 606
rect 882 605 883 606
rect 883 605 884 606
rect 885 605 886 606
rect 640 820 641 821
rect 642 820 643 821
rect 643 820 644 821
rect 645 820 646 821
rect 640 821 646 825
rect 640 825 641 826
rect 642 825 643 826
rect 643 825 644 826
rect 645 825 646 826
rect 720 720 721 721
rect 722 720 723 721
rect 723 720 724 721
rect 725 720 726 721
rect 720 721 726 725
rect 720 725 721 726
rect 722 725 723 726
rect 723 725 724 726
rect 725 725 726 726
rect 380 540 381 541
rect 382 540 383 541
rect 383 540 384 541
rect 385 540 386 541
rect 380 541 386 545
rect 380 545 381 546
rect 382 545 383 546
rect 383 545 384 546
rect 385 545 386 546
rect 440 600 441 601
rect 442 600 443 601
rect 443 600 444 601
rect 445 600 446 601
rect 440 601 446 605
rect 440 605 441 606
rect 442 605 443 606
rect 443 605 444 606
rect 445 605 446 606
rect 760 500 761 501
rect 762 500 763 501
rect 763 500 764 501
rect 765 500 766 501
rect 760 501 766 505
rect 760 505 761 506
rect 762 505 763 506
rect 763 505 764 506
rect 765 505 766 506
rect 600 420 601 421
rect 602 420 603 421
rect 603 420 604 421
rect 605 420 606 421
rect 600 421 606 425
rect 600 425 601 426
rect 602 425 603 426
rect 603 425 604 426
rect 605 425 606 426
rect 620 580 621 581
rect 622 580 623 581
rect 623 580 624 581
rect 625 580 626 581
rect 620 581 626 585
rect 620 585 621 586
rect 622 585 623 586
rect 623 585 624 586
rect 625 585 626 586
rect 700 360 701 361
rect 702 360 703 361
rect 703 360 704 361
rect 705 360 706 361
rect 700 361 706 365
rect 700 365 701 366
rect 702 365 703 366
rect 703 365 704 366
rect 705 365 706 366
rect 940 540 941 541
rect 942 540 943 541
rect 943 540 944 541
rect 945 540 946 541
rect 940 541 946 545
rect 940 545 941 546
rect 942 545 943 546
rect 943 545 944 546
rect 945 545 946 546
rect 340 760 341 761
rect 342 760 343 761
rect 343 760 344 761
rect 345 760 346 761
rect 340 761 346 765
rect 340 765 341 766
rect 342 765 343 766
rect 343 765 344 766
rect 345 765 346 766
rect 580 800 581 801
rect 582 800 583 801
rect 583 800 584 801
rect 585 800 586 801
rect 580 801 586 805
rect 580 805 581 806
rect 582 805 583 806
rect 583 805 584 806
rect 585 805 586 806
rect 500 660 501 661
rect 502 660 503 661
rect 503 660 504 661
rect 505 660 506 661
rect 500 661 506 665
rect 500 665 501 666
rect 502 665 503 666
rect 503 665 504 666
rect 505 665 506 666
rect 500 520 501 521
rect 502 520 503 521
rect 503 520 504 521
rect 505 520 506 521
rect 500 521 506 525
rect 500 525 501 526
rect 502 525 503 526
rect 503 525 504 526
rect 505 525 506 526
rect 660 320 661 321
rect 662 320 663 321
rect 663 320 664 321
rect 665 320 666 321
rect 660 321 666 325
rect 660 325 661 326
rect 662 325 663 326
rect 663 325 664 326
rect 665 325 666 326
rect 500 600 501 601
rect 502 600 503 601
rect 503 600 504 601
rect 505 600 506 601
rect 500 601 506 605
rect 500 605 501 606
rect 502 605 503 606
rect 503 605 504 606
rect 505 605 506 606
rect 660 420 661 421
rect 662 420 663 421
rect 663 420 664 421
rect 665 420 666 421
rect 660 421 666 425
rect 660 425 661 426
rect 662 425 663 426
rect 663 425 664 426
rect 665 425 666 426
rect 620 1060 621 1061
rect 622 1060 623 1061
rect 623 1060 624 1061
rect 625 1060 626 1061
rect 620 1061 626 1065
rect 620 1065 621 1066
rect 622 1065 623 1066
rect 623 1065 624 1066
rect 625 1065 626 1066
rect 520 520 521 521
rect 522 520 523 521
rect 523 520 524 521
rect 525 520 526 521
rect 520 521 526 525
rect 520 525 521 526
rect 522 525 523 526
rect 523 525 524 526
rect 525 525 526 526
rect 480 800 481 801
rect 482 800 483 801
rect 483 800 484 801
rect 485 800 486 801
rect 480 801 486 805
rect 480 805 481 806
rect 482 805 483 806
rect 483 805 484 806
rect 485 805 486 806
rect 460 540 461 541
rect 462 540 463 541
rect 463 540 464 541
rect 465 540 466 541
rect 460 541 466 545
rect 460 545 461 546
rect 462 545 463 546
rect 463 545 464 546
rect 465 545 466 546
rect 720 940 721 941
rect 722 940 723 941
rect 723 940 724 941
rect 725 940 726 941
rect 720 941 726 945
rect 720 945 721 946
rect 722 945 723 946
rect 723 945 724 946
rect 725 945 726 946
rect 900 580 901 581
rect 902 580 903 581
rect 903 580 904 581
rect 905 580 906 581
rect 900 581 906 585
rect 900 585 901 586
rect 902 585 903 586
rect 903 585 904 586
rect 905 585 906 586
rect 300 660 301 661
rect 302 660 303 661
rect 303 660 304 661
rect 305 660 306 661
rect 300 661 306 665
rect 300 665 301 666
rect 302 665 303 666
rect 303 665 304 666
rect 305 665 306 666
rect 520 420 521 421
rect 522 420 523 421
rect 523 420 524 421
rect 525 420 526 421
rect 520 421 526 425
rect 520 425 521 426
rect 522 425 523 426
rect 523 425 524 426
rect 525 425 526 426
rect 680 980 681 981
rect 682 980 683 981
rect 683 980 684 981
rect 685 980 686 981
rect 680 981 686 985
rect 680 985 681 986
rect 682 985 683 986
rect 683 985 684 986
rect 685 985 686 986
rect 420 680 421 681
rect 422 680 423 681
rect 423 680 424 681
rect 425 680 426 681
rect 420 681 426 685
rect 420 685 421 686
rect 422 685 423 686
rect 423 685 424 686
rect 425 685 426 686
rect 620 840 621 841
rect 622 840 623 841
rect 623 840 624 841
rect 625 840 626 841
rect 620 841 626 845
rect 620 845 621 846
rect 622 845 623 846
rect 623 845 624 846
rect 625 845 626 846
rect 980 700 981 701
rect 982 700 983 701
rect 983 700 984 701
rect 985 700 986 701
rect 980 701 986 705
rect 980 705 981 706
rect 982 705 983 706
rect 983 705 984 706
rect 985 705 986 706
rect 320 620 321 621
rect 322 620 323 621
rect 323 620 324 621
rect 325 620 326 621
rect 320 621 326 625
rect 320 625 321 626
rect 322 625 323 626
rect 323 625 324 626
rect 325 625 326 626
rect 380 640 381 641
rect 382 640 383 641
rect 383 640 384 641
rect 385 640 386 641
rect 380 641 386 645
rect 380 645 381 646
rect 382 645 383 646
rect 383 645 384 646
rect 385 645 386 646
rect 740 540 741 541
rect 742 540 743 541
rect 743 540 744 541
rect 745 540 746 541
rect 740 541 746 545
rect 740 545 741 546
rect 742 545 743 546
rect 743 545 744 546
rect 745 545 746 546
rect 400 620 401 621
rect 402 620 403 621
rect 403 620 404 621
rect 405 620 406 621
rect 400 621 406 625
rect 400 625 401 626
rect 402 625 403 626
rect 403 625 404 626
rect 405 625 406 626
rect 580 640 581 641
rect 582 640 583 641
rect 583 640 584 641
rect 585 640 586 641
rect 580 641 586 645
rect 580 645 581 646
rect 582 645 583 646
rect 583 645 584 646
rect 585 645 586 646
rect 620 1020 621 1021
rect 622 1020 623 1021
rect 623 1020 624 1021
rect 625 1020 626 1021
rect 620 1021 626 1025
rect 620 1025 621 1026
rect 622 1025 623 1026
rect 623 1025 624 1026
rect 625 1025 626 1026
rect 720 480 721 481
rect 722 480 723 481
rect 723 480 724 481
rect 725 480 726 481
rect 720 481 726 485
rect 720 485 721 486
rect 722 485 723 486
rect 723 485 724 486
rect 725 485 726 486
rect 340 580 341 581
rect 342 580 343 581
rect 343 580 344 581
rect 345 580 346 581
rect 340 581 346 585
rect 340 585 341 586
rect 342 585 343 586
rect 343 585 344 586
rect 345 585 346 586
rect 880 640 881 641
rect 882 640 883 641
rect 883 640 884 641
rect 885 640 886 641
rect 880 641 886 645
rect 880 645 881 646
rect 882 645 883 646
rect 883 645 884 646
rect 885 645 886 646
rect 580 400 581 401
rect 582 400 583 401
rect 583 400 584 401
rect 585 400 586 401
rect 580 401 586 405
rect 580 405 581 406
rect 582 405 583 406
rect 583 405 584 406
rect 585 405 586 406
rect 820 700 821 701
rect 822 700 823 701
rect 823 700 824 701
rect 825 700 826 701
rect 820 701 826 705
rect 820 705 821 706
rect 822 705 823 706
rect 823 705 824 706
rect 825 705 826 706
rect 500 760 501 761
rect 502 760 503 761
rect 503 760 504 761
rect 505 760 506 761
rect 500 761 506 765
rect 500 765 501 766
rect 502 765 503 766
rect 503 765 504 766
rect 505 765 506 766
rect 440 880 441 881
rect 442 880 443 881
rect 443 880 444 881
rect 445 880 446 881
rect 440 881 446 885
rect 440 885 441 886
rect 442 885 443 886
rect 443 885 444 886
rect 445 885 446 886
rect 760 440 761 441
rect 762 440 763 441
rect 763 440 764 441
rect 765 440 766 441
rect 760 441 766 445
rect 760 445 761 446
rect 762 445 763 446
rect 763 445 764 446
rect 765 445 766 446
rect 600 300 601 301
rect 602 300 603 301
rect 603 300 604 301
rect 605 300 606 301
rect 600 301 606 305
rect 600 305 601 306
rect 602 305 603 306
rect 603 305 604 306
rect 605 305 606 306
rect 960 700 961 701
rect 962 700 963 701
rect 963 700 964 701
rect 965 700 966 701
rect 960 701 966 705
rect 960 705 961 706
rect 962 705 963 706
rect 963 705 964 706
rect 965 705 966 706
rect 540 700 541 701
rect 542 700 543 701
rect 543 700 544 701
rect 545 700 546 701
rect 540 701 546 705
rect 540 705 541 706
rect 542 705 543 706
rect 543 705 544 706
rect 545 705 546 706
rect 840 900 841 901
rect 842 900 843 901
rect 843 900 844 901
rect 845 900 846 901
rect 840 901 846 905
rect 840 905 841 906
rect 842 905 843 906
rect 843 905 844 906
rect 845 905 846 906
rect 560 860 561 861
rect 562 860 563 861
rect 563 860 564 861
rect 565 860 566 861
rect 560 861 566 865
rect 560 865 561 866
rect 562 865 563 866
rect 563 865 564 866
rect 565 865 566 866
rect 680 440 681 441
rect 682 440 683 441
rect 683 440 684 441
rect 685 440 686 441
rect 680 441 686 445
rect 680 445 681 446
rect 682 445 683 446
rect 683 445 684 446
rect 685 445 686 446
rect 800 880 801 881
rect 802 880 803 881
rect 803 880 804 881
rect 805 880 806 881
rect 800 881 806 885
rect 800 885 801 886
rect 802 885 803 886
rect 803 885 804 886
rect 805 885 806 886
rect 780 520 781 521
rect 782 520 783 521
rect 783 520 784 521
rect 785 520 786 521
rect 780 521 786 525
rect 780 525 781 526
rect 782 525 783 526
rect 783 525 784 526
rect 785 525 786 526
rect 400 760 401 761
rect 402 760 403 761
rect 403 760 404 761
rect 405 760 406 761
rect 400 761 406 765
rect 400 765 401 766
rect 402 765 403 766
rect 403 765 404 766
rect 405 765 406 766
rect 720 280 721 281
rect 722 280 723 281
rect 723 280 724 281
rect 725 280 726 281
rect 720 281 726 285
rect 720 285 721 286
rect 722 285 723 286
rect 723 285 724 286
rect 725 285 726 286
rect 500 620 501 621
rect 502 620 503 621
rect 503 620 504 621
rect 505 620 506 621
rect 500 621 506 625
rect 500 625 501 626
rect 502 625 503 626
rect 503 625 504 626
rect 505 625 506 626
rect 460 500 461 501
rect 462 500 463 501
rect 463 500 464 501
rect 465 500 466 501
rect 460 501 466 505
rect 460 505 461 506
rect 462 505 463 506
rect 463 505 464 506
rect 465 505 466 506
rect 840 720 841 721
rect 842 720 843 721
rect 843 720 844 721
rect 845 720 846 721
rect 840 721 846 725
rect 840 725 841 726
rect 842 725 843 726
rect 843 725 844 726
rect 845 725 846 726
rect 620 1000 621 1001
rect 622 1000 623 1001
rect 623 1000 624 1001
rect 625 1000 626 1001
rect 620 1001 626 1005
rect 620 1005 621 1006
rect 622 1005 623 1006
rect 623 1005 624 1006
rect 625 1005 626 1006
rect 660 1000 661 1001
rect 662 1000 663 1001
rect 663 1000 664 1001
rect 665 1000 666 1001
rect 660 1001 666 1005
rect 660 1005 661 1006
rect 662 1005 663 1006
rect 663 1005 664 1006
rect 665 1005 666 1006
rect 560 640 561 641
rect 562 640 563 641
rect 563 640 564 641
rect 565 640 566 641
rect 560 641 566 645
rect 560 645 561 646
rect 562 645 563 646
rect 563 645 564 646
rect 565 645 566 646
rect 260 600 261 601
rect 262 600 263 601
rect 263 600 264 601
rect 265 600 266 601
rect 260 601 266 605
rect 260 605 261 606
rect 262 605 263 606
rect 263 605 264 606
rect 265 605 266 606
rect 400 560 401 561
rect 402 560 403 561
rect 403 560 404 561
rect 405 560 406 561
rect 400 561 406 565
rect 400 565 401 566
rect 402 565 403 566
rect 403 565 404 566
rect 405 565 406 566
rect 420 660 421 661
rect 422 660 423 661
rect 423 660 424 661
rect 425 660 426 661
rect 420 661 426 665
rect 420 665 421 666
rect 422 665 423 666
rect 423 665 424 666
rect 425 665 426 666
rect 260 660 261 661
rect 262 660 263 661
rect 263 660 264 661
rect 265 660 266 661
rect 260 661 266 665
rect 260 665 261 666
rect 262 665 263 666
rect 263 665 264 666
rect 265 665 266 666
rect 660 760 661 761
rect 662 760 663 761
rect 663 760 664 761
rect 665 760 666 761
rect 660 761 666 765
rect 660 765 661 766
rect 662 765 663 766
rect 663 765 664 766
rect 665 765 666 766
rect 1020 640 1021 641
rect 1022 640 1023 641
rect 1023 640 1024 641
rect 1025 640 1026 641
rect 1020 641 1026 645
rect 1020 645 1021 646
rect 1022 645 1023 646
rect 1023 645 1024 646
rect 1025 645 1026 646
rect 640 960 641 961
rect 642 960 643 961
rect 643 960 644 961
rect 645 960 646 961
rect 640 961 646 965
rect 640 965 641 966
rect 642 965 643 966
rect 643 965 644 966
rect 645 965 646 966
rect 300 760 301 761
rect 302 760 303 761
rect 303 760 304 761
rect 305 760 306 761
rect 300 761 306 765
rect 300 765 301 766
rect 302 765 303 766
rect 303 765 304 766
rect 305 765 306 766
rect 660 860 661 861
rect 662 860 663 861
rect 663 860 664 861
rect 665 860 666 861
rect 660 861 666 865
rect 660 865 661 866
rect 662 865 663 866
rect 663 865 664 866
rect 665 865 666 866
rect 960 540 961 541
rect 962 540 963 541
rect 963 540 964 541
rect 965 540 966 541
rect 960 541 966 545
rect 960 545 961 546
rect 962 545 963 546
rect 963 545 964 546
rect 965 545 966 546
rect 820 780 821 781
rect 822 780 823 781
rect 823 780 824 781
rect 825 780 826 781
rect 820 781 826 785
rect 820 785 821 786
rect 822 785 823 786
rect 823 785 824 786
rect 825 785 826 786
rect 840 880 841 881
rect 842 880 843 881
rect 843 880 844 881
rect 845 880 846 881
rect 840 881 846 885
rect 840 885 841 886
rect 842 885 843 886
rect 843 885 844 886
rect 845 885 846 886
rect 740 500 741 501
rect 742 500 743 501
rect 743 500 744 501
rect 745 500 746 501
rect 740 501 746 505
rect 740 505 741 506
rect 742 505 743 506
rect 743 505 744 506
rect 745 505 746 506
rect 620 420 621 421
rect 622 420 623 421
rect 623 420 624 421
rect 625 420 626 421
rect 620 421 626 425
rect 620 425 621 426
rect 622 425 623 426
rect 623 425 624 426
rect 625 425 626 426
rect 880 900 881 901
rect 882 900 883 901
rect 883 900 884 901
rect 885 900 886 901
rect 880 901 886 905
rect 880 905 881 906
rect 882 905 883 906
rect 883 905 884 906
rect 885 905 886 906
rect 280 620 281 621
rect 282 620 283 621
rect 283 620 284 621
rect 285 620 286 621
rect 280 621 286 625
rect 280 625 281 626
rect 282 625 283 626
rect 283 625 284 626
rect 285 625 286 626
rect 640 340 641 341
rect 642 340 643 341
rect 643 340 644 341
rect 645 340 646 341
rect 640 341 646 345
rect 640 345 641 346
rect 642 345 643 346
rect 643 345 644 346
rect 645 345 646 346
rect 540 620 541 621
rect 542 620 543 621
rect 543 620 544 621
rect 545 620 546 621
rect 540 621 546 625
rect 540 625 541 626
rect 542 625 543 626
rect 543 625 544 626
rect 545 625 546 626
rect 480 620 481 621
rect 482 620 483 621
rect 483 620 484 621
rect 485 620 486 621
rect 480 621 486 625
rect 480 625 481 626
rect 482 625 483 626
rect 483 625 484 626
rect 485 625 486 626
rect 480 420 481 421
rect 482 420 483 421
rect 483 420 484 421
rect 485 420 486 421
rect 480 421 486 425
rect 480 425 481 426
rect 482 425 483 426
rect 483 425 484 426
rect 485 425 486 426
rect 240 680 241 681
rect 242 680 243 681
rect 243 680 244 681
rect 245 680 246 681
rect 240 681 246 685
rect 240 685 241 686
rect 242 685 243 686
rect 243 685 244 686
rect 245 685 246 686
rect 600 820 601 821
rect 602 820 603 821
rect 603 820 604 821
rect 605 820 606 821
rect 600 821 606 825
rect 600 825 601 826
rect 602 825 603 826
rect 603 825 604 826
rect 605 825 606 826
rect 560 620 561 621
rect 562 620 563 621
rect 563 620 564 621
rect 565 620 566 621
rect 560 621 566 625
rect 560 625 561 626
rect 562 625 563 626
rect 563 625 564 626
rect 565 625 566 626
rect 900 820 901 821
rect 902 820 903 821
rect 903 820 904 821
rect 905 820 906 821
rect 900 821 906 825
rect 900 825 901 826
rect 902 825 903 826
rect 903 825 904 826
rect 905 825 906 826
rect 800 940 801 941
rect 802 940 803 941
rect 803 940 804 941
rect 805 940 806 941
rect 800 941 806 945
rect 800 945 801 946
rect 802 945 803 946
rect 803 945 804 946
rect 805 945 806 946
rect 820 480 821 481
rect 822 480 823 481
rect 823 480 824 481
rect 825 480 826 481
rect 820 481 826 485
rect 820 485 821 486
rect 822 485 823 486
rect 823 485 824 486
rect 825 485 826 486
rect 1000 700 1001 701
rect 1002 700 1003 701
rect 1003 700 1004 701
rect 1005 700 1006 701
rect 1000 701 1006 705
rect 1000 705 1001 706
rect 1002 705 1003 706
rect 1003 705 1004 706
rect 1005 705 1006 706
rect 320 680 321 681
rect 322 680 323 681
rect 323 680 324 681
rect 325 680 326 681
rect 320 681 326 685
rect 320 685 321 686
rect 322 685 323 686
rect 323 685 324 686
rect 325 685 326 686
rect 740 380 741 381
rect 742 380 743 381
rect 743 380 744 381
rect 745 380 746 381
rect 740 381 746 385
rect 740 385 741 386
rect 742 385 743 386
rect 743 385 744 386
rect 745 385 746 386
rect 940 820 941 821
rect 942 820 943 821
rect 943 820 944 821
rect 945 820 946 821
rect 940 821 946 825
rect 940 825 941 826
rect 942 825 943 826
rect 943 825 944 826
rect 945 825 946 826
rect 740 1040 741 1041
rect 742 1040 743 1041
rect 743 1040 744 1041
rect 745 1040 746 1041
rect 740 1041 746 1045
rect 740 1045 741 1046
rect 742 1045 743 1046
rect 743 1045 744 1046
rect 745 1045 746 1046
rect 420 520 421 521
rect 422 520 423 521
rect 423 520 424 521
rect 425 520 426 521
rect 420 521 426 525
rect 420 525 421 526
rect 422 525 423 526
rect 423 525 424 526
rect 425 525 426 526
rect 780 940 781 941
rect 782 940 783 941
rect 783 940 784 941
rect 785 940 786 941
rect 780 941 786 945
rect 780 945 781 946
rect 782 945 783 946
rect 783 945 784 946
rect 785 945 786 946
rect 900 480 901 481
rect 902 480 903 481
rect 903 480 904 481
rect 905 480 906 481
rect 900 481 906 485
rect 900 485 901 486
rect 902 485 903 486
rect 903 485 904 486
rect 905 485 906 486
rect 740 400 741 401
rect 742 400 743 401
rect 743 400 744 401
rect 745 400 746 401
rect 740 401 746 405
rect 740 405 741 406
rect 742 405 743 406
rect 743 405 744 406
rect 745 405 746 406
rect 880 760 881 761
rect 882 760 883 761
rect 883 760 884 761
rect 885 760 886 761
rect 880 761 886 765
rect 880 765 881 766
rect 882 765 883 766
rect 883 765 884 766
rect 885 765 886 766
rect 700 1000 701 1001
rect 702 1000 703 1001
rect 703 1000 704 1001
rect 705 1000 706 1001
rect 700 1001 706 1005
rect 700 1005 701 1006
rect 702 1005 703 1006
rect 703 1005 704 1006
rect 705 1005 706 1006
rect 640 560 641 561
rect 642 560 643 561
rect 643 560 644 561
rect 645 560 646 561
rect 640 561 646 565
rect 640 565 641 566
rect 642 565 643 566
rect 643 565 644 566
rect 645 565 646 566
rect 600 320 601 321
rect 602 320 603 321
rect 603 320 604 321
rect 605 320 606 321
rect 600 321 606 325
rect 600 325 601 326
rect 602 325 603 326
rect 603 325 604 326
rect 605 325 606 326
rect 760 380 761 381
rect 762 380 763 381
rect 763 380 764 381
rect 765 380 766 381
rect 760 381 766 385
rect 760 385 761 386
rect 762 385 763 386
rect 763 385 764 386
rect 765 385 766 386
rect 840 500 841 501
rect 842 500 843 501
rect 843 500 844 501
rect 845 500 846 501
rect 840 501 846 505
rect 840 505 841 506
rect 842 505 843 506
rect 843 505 844 506
rect 845 505 846 506
rect 940 560 941 561
rect 942 560 943 561
rect 943 560 944 561
rect 945 560 946 561
rect 940 561 946 565
rect 940 565 941 566
rect 942 565 943 566
rect 943 565 944 566
rect 945 565 946 566
rect 1060 660 1061 661
rect 1062 660 1063 661
rect 1063 660 1064 661
rect 1065 660 1066 661
rect 1060 661 1066 665
rect 1060 665 1061 666
rect 1062 665 1063 666
rect 1063 665 1064 666
rect 1065 665 1066 666
rect 600 720 601 721
rect 602 720 603 721
rect 603 720 604 721
rect 605 720 606 721
rect 600 721 606 725
rect 600 725 601 726
rect 602 725 603 726
rect 603 725 604 726
rect 605 725 606 726
rect 440 520 441 521
rect 442 520 443 521
rect 443 520 444 521
rect 445 520 446 521
rect 440 521 446 525
rect 440 525 441 526
rect 442 525 443 526
rect 443 525 444 526
rect 445 525 446 526
rect 740 760 741 761
rect 742 760 743 761
rect 743 760 744 761
rect 745 760 746 761
rect 740 761 746 765
rect 740 765 741 766
rect 742 765 743 766
rect 743 765 744 766
rect 745 765 746 766
rect 340 560 341 561
rect 342 560 343 561
rect 343 560 344 561
rect 345 560 346 561
rect 340 561 346 565
rect 340 565 341 566
rect 342 565 343 566
rect 343 565 344 566
rect 345 565 346 566
rect 360 560 361 561
rect 362 560 363 561
rect 363 560 364 561
rect 365 560 366 561
rect 360 561 366 565
rect 360 565 361 566
rect 362 565 363 566
rect 363 565 364 566
rect 365 565 366 566
rect 820 400 821 401
rect 822 400 823 401
rect 823 400 824 401
rect 825 400 826 401
rect 820 401 826 405
rect 820 405 821 406
rect 822 405 823 406
rect 823 405 824 406
rect 825 405 826 406
rect 640 1080 641 1081
rect 642 1080 643 1081
rect 643 1080 644 1081
rect 645 1080 646 1081
rect 640 1081 646 1085
rect 640 1085 641 1086
rect 642 1085 643 1086
rect 643 1085 644 1086
rect 645 1085 646 1086
rect 680 520 681 521
rect 682 520 683 521
rect 683 520 684 521
rect 685 520 686 521
rect 680 521 686 525
rect 680 525 681 526
rect 682 525 683 526
rect 683 525 684 526
rect 685 525 686 526
rect 760 640 761 641
rect 762 640 763 641
rect 763 640 764 641
rect 765 640 766 641
rect 760 641 766 645
rect 760 645 761 646
rect 762 645 763 646
rect 763 645 764 646
rect 765 645 766 646
rect 820 820 821 821
rect 822 820 823 821
rect 823 820 824 821
rect 825 820 826 821
rect 820 821 826 825
rect 820 825 821 826
rect 822 825 823 826
rect 823 825 824 826
rect 825 825 826 826
rect 760 420 761 421
rect 762 420 763 421
rect 763 420 764 421
rect 765 420 766 421
rect 760 421 766 425
rect 760 425 761 426
rect 762 425 763 426
rect 763 425 764 426
rect 765 425 766 426
rect 500 880 501 881
rect 502 880 503 881
rect 503 880 504 881
rect 505 880 506 881
rect 500 881 506 885
rect 500 885 501 886
rect 502 885 503 886
rect 503 885 504 886
rect 505 885 506 886
rect 620 600 621 601
rect 622 600 623 601
rect 623 600 624 601
rect 625 600 626 601
rect 620 601 626 605
rect 620 605 621 606
rect 622 605 623 606
rect 623 605 624 606
rect 625 605 626 606
rect 260 700 261 701
rect 262 700 263 701
rect 263 700 264 701
rect 265 700 266 701
rect 260 701 266 705
rect 260 705 261 706
rect 262 705 263 706
rect 263 705 264 706
rect 265 705 266 706
rect 800 500 801 501
rect 802 500 803 501
rect 803 500 804 501
rect 805 500 806 501
rect 800 501 806 505
rect 800 505 801 506
rect 802 505 803 506
rect 803 505 804 506
rect 805 505 806 506
rect 420 800 421 801
rect 422 800 423 801
rect 423 800 424 801
rect 425 800 426 801
rect 420 801 426 805
rect 420 805 421 806
rect 422 805 423 806
rect 423 805 424 806
rect 425 805 426 806
rect 860 440 861 441
rect 862 440 863 441
rect 863 440 864 441
rect 865 440 866 441
rect 860 441 866 445
rect 860 445 861 446
rect 862 445 863 446
rect 863 445 864 446
rect 865 445 866 446
rect 760 1040 761 1041
rect 762 1040 763 1041
rect 763 1040 764 1041
rect 765 1040 766 1041
rect 760 1041 766 1045
rect 760 1045 761 1046
rect 762 1045 763 1046
rect 763 1045 764 1046
rect 765 1045 766 1046
rect 820 920 821 921
rect 822 920 823 921
rect 823 920 824 921
rect 825 920 826 921
rect 820 921 826 925
rect 820 925 821 926
rect 822 925 823 926
rect 823 925 824 926
rect 825 925 826 926
rect 680 780 681 781
rect 682 780 683 781
rect 683 780 684 781
rect 685 780 686 781
rect 680 781 686 785
rect 680 785 681 786
rect 682 785 683 786
rect 683 785 684 786
rect 685 785 686 786
rect 660 500 661 501
rect 662 500 663 501
rect 663 500 664 501
rect 665 500 666 501
rect 660 501 666 505
rect 660 505 661 506
rect 662 505 663 506
rect 663 505 664 506
rect 665 505 666 506
rect 720 980 721 981
rect 722 980 723 981
rect 723 980 724 981
rect 725 980 726 981
rect 720 981 726 985
rect 720 985 721 986
rect 722 985 723 986
rect 723 985 724 986
rect 725 985 726 986
rect 580 660 581 661
rect 582 660 583 661
rect 583 660 584 661
rect 585 660 586 661
rect 580 661 586 665
rect 580 665 581 666
rect 582 665 583 666
rect 583 665 584 666
rect 585 665 586 666
rect 940 760 941 761
rect 942 760 943 761
rect 943 760 944 761
rect 945 760 946 761
rect 940 761 946 765
rect 940 765 941 766
rect 942 765 943 766
rect 943 765 944 766
rect 945 765 946 766
rect 860 540 861 541
rect 862 540 863 541
rect 863 540 864 541
rect 865 540 866 541
rect 860 541 866 545
rect 860 545 861 546
rect 862 545 863 546
rect 863 545 864 546
rect 865 545 866 546
rect 1040 640 1041 641
rect 1042 640 1043 641
rect 1043 640 1044 641
rect 1045 640 1046 641
rect 1040 641 1046 645
rect 1040 645 1041 646
rect 1042 645 1043 646
rect 1043 645 1044 646
rect 1045 645 1046 646
rect 700 820 701 821
rect 702 820 703 821
rect 703 820 704 821
rect 705 820 706 821
rect 700 821 706 825
rect 700 825 701 826
rect 702 825 703 826
rect 703 825 704 826
rect 705 825 706 826
rect 820 860 821 861
rect 822 860 823 861
rect 823 860 824 861
rect 825 860 826 861
rect 820 861 826 865
rect 820 865 821 866
rect 822 865 823 866
rect 823 865 824 866
rect 825 865 826 866
rect 960 620 961 621
rect 962 620 963 621
rect 963 620 964 621
rect 965 620 966 621
rect 960 621 966 625
rect 960 625 961 626
rect 962 625 963 626
rect 963 625 964 626
rect 965 625 966 626
rect 540 380 541 381
rect 542 380 543 381
rect 543 380 544 381
rect 545 380 546 381
rect 540 381 546 385
rect 540 385 541 386
rect 542 385 543 386
rect 543 385 544 386
rect 545 385 546 386
rect 700 940 701 941
rect 702 940 703 941
rect 703 940 704 941
rect 705 940 706 941
rect 700 941 706 945
rect 700 945 701 946
rect 702 945 703 946
rect 703 945 704 946
rect 705 945 706 946
rect 640 660 641 661
rect 642 660 643 661
rect 643 660 644 661
rect 645 660 646 661
rect 640 661 646 665
rect 640 665 641 666
rect 642 665 643 666
rect 643 665 644 666
rect 645 665 646 666
rect 700 880 701 881
rect 702 880 703 881
rect 703 880 704 881
rect 705 880 706 881
rect 700 881 706 885
rect 700 885 701 886
rect 702 885 703 886
rect 703 885 704 886
rect 705 885 706 886
rect 660 540 661 541
rect 662 540 663 541
rect 663 540 664 541
rect 665 540 666 541
rect 660 541 666 545
rect 660 545 661 546
rect 662 545 663 546
rect 663 545 664 546
rect 665 545 666 546
rect 740 680 741 681
rect 742 680 743 681
rect 743 680 744 681
rect 745 680 746 681
rect 740 681 746 685
rect 740 685 741 686
rect 742 685 743 686
rect 743 685 744 686
rect 745 685 746 686
rect 620 340 621 341
rect 622 340 623 341
rect 623 340 624 341
rect 625 340 626 341
rect 620 341 626 345
rect 620 345 621 346
rect 622 345 623 346
rect 623 345 624 346
rect 625 345 626 346
rect 880 580 881 581
rect 882 580 883 581
rect 883 580 884 581
rect 885 580 886 581
rect 880 581 886 585
rect 880 585 881 586
rect 882 585 883 586
rect 883 585 884 586
rect 885 585 886 586
rect 700 760 701 761
rect 702 760 703 761
rect 703 760 704 761
rect 705 760 706 761
rect 700 761 706 765
rect 700 765 701 766
rect 702 765 703 766
rect 703 765 704 766
rect 705 765 706 766
rect 700 720 701 721
rect 702 720 703 721
rect 703 720 704 721
rect 705 720 706 721
rect 700 721 706 725
rect 700 725 701 726
rect 702 725 703 726
rect 703 725 704 726
rect 705 725 706 726
rect 600 560 601 561
rect 602 560 603 561
rect 603 560 604 561
rect 605 560 606 561
rect 600 561 606 565
rect 600 565 601 566
rect 602 565 603 566
rect 603 565 604 566
rect 605 565 606 566
rect 580 1040 581 1041
rect 582 1040 583 1041
rect 583 1040 584 1041
rect 585 1040 586 1041
rect 580 1041 586 1045
rect 580 1045 581 1046
rect 582 1045 583 1046
rect 583 1045 584 1046
rect 585 1045 586 1046
rect 720 540 721 541
rect 722 540 723 541
rect 723 540 724 541
rect 725 540 726 541
rect 720 541 726 545
rect 720 545 721 546
rect 722 545 723 546
rect 723 545 724 546
rect 725 545 726 546
rect 620 520 621 521
rect 622 520 623 521
rect 623 520 624 521
rect 625 520 626 521
rect 620 521 626 525
rect 620 525 621 526
rect 622 525 623 526
rect 623 525 624 526
rect 625 525 626 526
rect 640 780 641 781
rect 642 780 643 781
rect 643 780 644 781
rect 645 780 646 781
rect 640 781 646 785
rect 640 785 641 786
rect 642 785 643 786
rect 643 785 644 786
rect 645 785 646 786
rect 520 580 521 581
rect 522 580 523 581
rect 523 580 524 581
rect 525 580 526 581
rect 520 581 526 585
rect 520 585 521 586
rect 522 585 523 586
rect 523 585 524 586
rect 525 585 526 586
rect 520 660 521 661
rect 522 660 523 661
rect 523 660 524 661
rect 525 660 526 661
rect 520 661 526 665
rect 520 665 521 666
rect 522 665 523 666
rect 523 665 524 666
rect 525 665 526 666
rect 800 860 801 861
rect 802 860 803 861
rect 803 860 804 861
rect 805 860 806 861
rect 800 861 806 865
rect 800 865 801 866
rect 802 865 803 866
rect 803 865 804 866
rect 805 865 806 866
rect 320 600 321 601
rect 322 600 323 601
rect 323 600 324 601
rect 325 600 326 601
rect 320 601 326 605
rect 320 605 321 606
rect 322 605 323 606
rect 323 605 324 606
rect 325 605 326 606
rect 540 460 541 461
rect 542 460 543 461
rect 543 460 544 461
rect 545 460 546 461
rect 540 461 546 465
rect 540 465 541 466
rect 542 465 543 466
rect 543 465 544 466
rect 545 465 546 466
rect 800 900 801 901
rect 802 900 803 901
rect 803 900 804 901
rect 805 900 806 901
rect 800 901 806 905
rect 800 905 801 906
rect 802 905 803 906
rect 803 905 804 906
rect 805 905 806 906
rect 600 1000 601 1001
rect 602 1000 603 1001
rect 603 1000 604 1001
rect 605 1000 606 1001
rect 600 1001 606 1005
rect 600 1005 601 1006
rect 602 1005 603 1006
rect 603 1005 604 1006
rect 605 1005 606 1006
rect 440 860 441 861
rect 442 860 443 861
rect 443 860 444 861
rect 445 860 446 861
rect 440 861 446 865
rect 440 865 441 866
rect 442 865 443 866
rect 443 865 444 866
rect 445 865 446 866
rect 720 420 721 421
rect 722 420 723 421
rect 723 420 724 421
rect 725 420 726 421
rect 720 421 726 425
rect 720 425 721 426
rect 722 425 723 426
rect 723 425 724 426
rect 725 425 726 426
rect 580 720 581 721
rect 582 720 583 721
rect 583 720 584 721
rect 585 720 586 721
rect 580 721 586 725
rect 580 725 581 726
rect 582 725 583 726
rect 583 725 584 726
rect 585 725 586 726
rect 740 660 741 661
rect 742 660 743 661
rect 743 660 744 661
rect 745 660 746 661
rect 740 661 746 665
rect 740 665 741 666
rect 742 665 743 666
rect 743 665 744 666
rect 745 665 746 666
rect 820 620 821 621
rect 822 620 823 621
rect 823 620 824 621
rect 825 620 826 621
rect 820 621 826 625
rect 820 625 821 626
rect 822 625 823 626
rect 823 625 824 626
rect 825 625 826 626
rect 360 720 361 721
rect 362 720 363 721
rect 363 720 364 721
rect 365 720 366 721
rect 360 721 366 725
rect 360 725 361 726
rect 362 725 363 726
rect 363 725 364 726
rect 365 725 366 726
rect 540 940 541 941
rect 542 940 543 941
rect 543 940 544 941
rect 545 940 546 941
rect 540 941 546 945
rect 540 945 541 946
rect 542 945 543 946
rect 543 945 544 946
rect 545 945 546 946
rect 540 680 541 681
rect 542 680 543 681
rect 543 680 544 681
rect 545 680 546 681
rect 540 681 546 685
rect 540 685 541 686
rect 542 685 543 686
rect 543 685 544 686
rect 545 685 546 686
rect 960 640 961 641
rect 962 640 963 641
rect 963 640 964 641
rect 965 640 966 641
rect 960 641 966 645
rect 960 645 961 646
rect 962 645 963 646
rect 963 645 964 646
rect 965 645 966 646
rect 580 840 581 841
rect 582 840 583 841
rect 583 840 584 841
rect 585 840 586 841
rect 580 841 586 845
rect 580 845 581 846
rect 582 845 583 846
rect 583 845 584 846
rect 585 845 586 846
rect 720 900 721 901
rect 722 900 723 901
rect 723 900 724 901
rect 725 900 726 901
rect 720 901 726 905
rect 720 905 721 906
rect 722 905 723 906
rect 723 905 724 906
rect 725 905 726 906
rect 660 840 661 841
rect 662 840 663 841
rect 663 840 664 841
rect 665 840 666 841
rect 660 841 666 845
rect 660 845 661 846
rect 662 845 663 846
rect 663 845 664 846
rect 665 845 666 846
rect 700 300 701 301
rect 702 300 703 301
rect 703 300 704 301
rect 705 300 706 301
rect 700 301 706 305
rect 700 305 701 306
rect 702 305 703 306
rect 703 305 704 306
rect 705 305 706 306
rect 440 760 441 761
rect 442 760 443 761
rect 443 760 444 761
rect 445 760 446 761
rect 440 761 446 765
rect 440 765 441 766
rect 442 765 443 766
rect 443 765 444 766
rect 445 765 446 766
rect 440 540 441 541
rect 442 540 443 541
rect 443 540 444 541
rect 445 540 446 541
rect 440 541 446 545
rect 440 545 441 546
rect 442 545 443 546
rect 443 545 444 546
rect 445 545 446 546
rect 460 460 461 461
rect 462 460 463 461
rect 463 460 464 461
rect 465 460 466 461
rect 460 461 466 465
rect 460 465 461 466
rect 462 465 463 466
rect 463 465 464 466
rect 465 465 466 466
rect 400 700 401 701
rect 402 700 403 701
rect 403 700 404 701
rect 405 700 406 701
rect 400 701 406 705
rect 400 705 401 706
rect 402 705 403 706
rect 403 705 404 706
rect 405 705 406 706
rect 680 480 681 481
rect 682 480 683 481
rect 683 480 684 481
rect 685 480 686 481
rect 680 481 686 485
rect 680 485 681 486
rect 682 485 683 486
rect 683 485 684 486
rect 685 485 686 486
rect 680 340 681 341
rect 682 340 683 341
rect 683 340 684 341
rect 685 340 686 341
rect 680 341 686 345
rect 680 345 681 346
rect 682 345 683 346
rect 683 345 684 346
rect 685 345 686 346
rect 720 920 721 921
rect 722 920 723 921
rect 723 920 724 921
rect 725 920 726 921
rect 720 921 726 925
rect 720 925 721 926
rect 722 925 723 926
rect 723 925 724 926
rect 725 925 726 926
rect 540 860 541 861
rect 542 860 543 861
rect 543 860 544 861
rect 545 860 546 861
rect 540 861 546 865
rect 540 865 541 866
rect 542 865 543 866
rect 543 865 544 866
rect 545 865 546 866
rect 700 1040 701 1041
rect 702 1040 703 1041
rect 703 1040 704 1041
rect 705 1040 706 1041
rect 700 1041 706 1045
rect 700 1045 701 1046
rect 702 1045 703 1046
rect 703 1045 704 1046
rect 705 1045 706 1046
rect 780 980 781 981
rect 782 980 783 981
rect 783 980 784 981
rect 785 980 786 981
rect 780 981 786 985
rect 780 985 781 986
rect 782 985 783 986
rect 783 985 784 986
rect 785 985 786 986
rect 920 520 921 521
rect 922 520 923 521
rect 923 520 924 521
rect 925 520 926 521
rect 920 521 926 525
rect 920 525 921 526
rect 922 525 923 526
rect 923 525 924 526
rect 925 525 926 526
rect 460 600 461 601
rect 462 600 463 601
rect 463 600 464 601
rect 465 600 466 601
rect 460 601 466 605
rect 460 605 461 606
rect 462 605 463 606
rect 463 605 464 606
rect 465 605 466 606
rect 860 680 861 681
rect 862 680 863 681
rect 863 680 864 681
rect 865 680 866 681
rect 860 681 866 685
rect 860 685 861 686
rect 862 685 863 686
rect 863 685 864 686
rect 865 685 866 686
rect 660 740 661 741
rect 662 740 663 741
rect 663 740 664 741
rect 665 740 666 741
rect 660 741 666 745
rect 660 745 661 746
rect 662 745 663 746
rect 663 745 664 746
rect 665 745 666 746
rect 480 580 481 581
rect 482 580 483 581
rect 483 580 484 581
rect 485 580 486 581
rect 480 581 486 585
rect 480 585 481 586
rect 482 585 483 586
rect 483 585 484 586
rect 485 585 486 586
rect 820 640 821 641
rect 822 640 823 641
rect 823 640 824 641
rect 825 640 826 641
rect 820 641 826 645
rect 820 645 821 646
rect 822 645 823 646
rect 823 645 824 646
rect 825 645 826 646
rect 320 740 321 741
rect 322 740 323 741
rect 323 740 324 741
rect 325 740 326 741
rect 320 741 326 745
rect 320 745 321 746
rect 322 745 323 746
rect 323 745 324 746
rect 325 745 326 746
rect 640 900 641 901
rect 642 900 643 901
rect 643 900 644 901
rect 645 900 646 901
rect 640 901 646 905
rect 640 905 641 906
rect 642 905 643 906
rect 643 905 644 906
rect 645 905 646 906
rect 660 960 661 961
rect 662 960 663 961
rect 663 960 664 961
rect 665 960 666 961
rect 660 961 666 965
rect 660 965 661 966
rect 662 965 663 966
rect 663 965 664 966
rect 665 965 666 966
rect 600 540 601 541
rect 602 540 603 541
rect 603 540 604 541
rect 605 540 606 541
rect 600 541 606 545
rect 600 545 601 546
rect 602 545 603 546
rect 603 545 604 546
rect 605 545 606 546
rect 440 460 441 461
rect 442 460 443 461
rect 443 460 444 461
rect 445 460 446 461
rect 440 461 446 465
rect 440 465 441 466
rect 442 465 443 466
rect 443 465 444 466
rect 445 465 446 466
rect 680 360 681 361
rect 682 360 683 361
rect 683 360 684 361
rect 685 360 686 361
rect 680 361 686 365
rect 680 365 681 366
rect 682 365 683 366
rect 683 365 684 366
rect 685 365 686 366
rect 820 660 821 661
rect 822 660 823 661
rect 823 660 824 661
rect 825 660 826 661
rect 820 661 826 665
rect 820 665 821 666
rect 822 665 823 666
rect 823 665 824 666
rect 825 665 826 666
rect 740 860 741 861
rect 742 860 743 861
rect 743 860 744 861
rect 745 860 746 861
rect 740 861 746 865
rect 740 865 741 866
rect 742 865 743 866
rect 743 865 744 866
rect 745 865 746 866
rect 620 300 621 301
rect 622 300 623 301
rect 623 300 624 301
rect 625 300 626 301
rect 620 301 626 305
rect 620 305 621 306
rect 622 305 623 306
rect 623 305 624 306
rect 625 305 626 306
rect 740 580 741 581
rect 742 580 743 581
rect 743 580 744 581
rect 745 580 746 581
rect 740 581 746 585
rect 740 585 741 586
rect 742 585 743 586
rect 743 585 744 586
rect 745 585 746 586
rect 840 660 841 661
rect 842 660 843 661
rect 843 660 844 661
rect 845 660 846 661
rect 840 661 846 665
rect 840 665 841 666
rect 842 665 843 666
rect 843 665 844 666
rect 845 665 846 666
rect 240 640 241 641
rect 242 640 243 641
rect 243 640 244 641
rect 245 640 246 641
rect 240 641 246 645
rect 240 645 241 646
rect 242 645 243 646
rect 243 645 244 646
rect 245 645 246 646
rect 800 600 801 601
rect 802 600 803 601
rect 803 600 804 601
rect 805 600 806 601
rect 800 601 806 605
rect 800 605 801 606
rect 802 605 803 606
rect 803 605 804 606
rect 805 605 806 606
rect 740 740 741 741
rect 742 740 743 741
rect 743 740 744 741
rect 745 740 746 741
rect 740 741 746 745
rect 740 745 741 746
rect 742 745 743 746
rect 743 745 744 746
rect 745 745 746 746
rect 680 540 681 541
rect 682 540 683 541
rect 683 540 684 541
rect 685 540 686 541
rect 680 541 686 545
rect 680 545 681 546
rect 682 545 683 546
rect 683 545 684 546
rect 685 545 686 546
rect 980 720 981 721
rect 982 720 983 721
rect 983 720 984 721
rect 985 720 986 721
rect 980 721 986 725
rect 980 725 981 726
rect 982 725 983 726
rect 983 725 984 726
rect 985 725 986 726
rect 1020 740 1021 741
rect 1022 740 1023 741
rect 1023 740 1024 741
rect 1025 740 1026 741
rect 1020 741 1026 745
rect 1020 745 1021 746
rect 1022 745 1023 746
rect 1023 745 1024 746
rect 1025 745 1026 746
rect 460 420 461 421
rect 462 420 463 421
rect 463 420 464 421
rect 465 420 466 421
rect 460 421 466 425
rect 460 425 461 426
rect 462 425 463 426
rect 463 425 464 426
rect 465 425 466 426
rect 500 400 501 401
rect 502 400 503 401
rect 503 400 504 401
rect 505 400 506 401
rect 500 401 506 405
rect 500 405 501 406
rect 502 405 503 406
rect 503 405 504 406
rect 505 405 506 406
rect 400 720 401 721
rect 402 720 403 721
rect 403 720 404 721
rect 405 720 406 721
rect 400 721 406 725
rect 400 725 401 726
rect 402 725 403 726
rect 403 725 404 726
rect 405 725 406 726
rect 940 840 941 841
rect 942 840 943 841
rect 943 840 944 841
rect 945 840 946 841
rect 940 841 946 845
rect 940 845 941 846
rect 942 845 943 846
rect 943 845 944 846
rect 945 845 946 846
rect 720 380 721 381
rect 722 380 723 381
rect 723 380 724 381
rect 725 380 726 381
rect 720 381 726 385
rect 720 385 721 386
rect 722 385 723 386
rect 723 385 724 386
rect 725 385 726 386
rect 300 620 301 621
rect 302 620 303 621
rect 303 620 304 621
rect 305 620 306 621
rect 300 621 306 625
rect 300 625 301 626
rect 302 625 303 626
rect 303 625 304 626
rect 305 625 306 626
rect 700 420 701 421
rect 702 420 703 421
rect 703 420 704 421
rect 705 420 706 421
rect 700 421 706 425
rect 700 425 701 426
rect 702 425 703 426
rect 703 425 704 426
rect 705 425 706 426
rect 520 800 521 801
rect 522 800 523 801
rect 523 800 524 801
rect 525 800 526 801
rect 520 801 526 805
rect 520 805 521 806
rect 522 805 523 806
rect 523 805 524 806
rect 525 805 526 806
rect 520 480 521 481
rect 522 480 523 481
rect 523 480 524 481
rect 525 480 526 481
rect 520 481 526 485
rect 520 485 521 486
rect 522 485 523 486
rect 523 485 524 486
rect 525 485 526 486
rect 1000 640 1001 641
rect 1002 640 1003 641
rect 1003 640 1004 641
rect 1005 640 1006 641
rect 1000 641 1006 645
rect 1000 645 1001 646
rect 1002 645 1003 646
rect 1003 645 1004 646
rect 1005 645 1006 646
rect 460 580 461 581
rect 462 580 463 581
rect 463 580 464 581
rect 465 580 466 581
rect 460 581 466 585
rect 460 585 461 586
rect 462 585 463 586
rect 463 585 464 586
rect 465 585 466 586
rect 620 700 621 701
rect 622 700 623 701
rect 623 700 624 701
rect 625 700 626 701
rect 620 701 626 705
rect 620 705 621 706
rect 622 705 623 706
rect 623 705 624 706
rect 625 705 626 706
rect 920 740 921 741
rect 922 740 923 741
rect 923 740 924 741
rect 925 740 926 741
rect 920 741 926 745
rect 920 745 921 746
rect 922 745 923 746
rect 923 745 924 746
rect 925 745 926 746
rect 560 440 561 441
rect 562 440 563 441
rect 563 440 564 441
rect 565 440 566 441
rect 560 441 566 445
rect 560 445 561 446
rect 562 445 563 446
rect 563 445 564 446
rect 565 445 566 446
rect 640 1040 641 1041
rect 642 1040 643 1041
rect 643 1040 644 1041
rect 645 1040 646 1041
rect 640 1041 646 1045
rect 640 1045 641 1046
rect 642 1045 643 1046
rect 643 1045 644 1046
rect 645 1045 646 1046
rect 840 420 841 421
rect 842 420 843 421
rect 843 420 844 421
rect 845 420 846 421
rect 840 421 846 425
rect 840 425 841 426
rect 842 425 843 426
rect 843 425 844 426
rect 845 425 846 426
rect 420 820 421 821
rect 422 820 423 821
rect 423 820 424 821
rect 425 820 426 821
rect 420 821 426 825
rect 420 825 421 826
rect 422 825 423 826
rect 423 825 424 826
rect 425 825 426 826
rect 840 700 841 701
rect 842 700 843 701
rect 843 700 844 701
rect 845 700 846 701
rect 840 701 846 705
rect 840 705 841 706
rect 842 705 843 706
rect 843 705 844 706
rect 845 705 846 706
rect 600 780 601 781
rect 602 780 603 781
rect 603 780 604 781
rect 605 780 606 781
rect 600 781 606 785
rect 600 785 601 786
rect 602 785 603 786
rect 603 785 604 786
rect 605 785 606 786
rect 1060 700 1061 701
rect 1062 700 1063 701
rect 1063 700 1064 701
rect 1065 700 1066 701
rect 1060 701 1066 705
rect 1060 705 1061 706
rect 1062 705 1063 706
rect 1063 705 1064 706
rect 1065 705 1066 706
rect 720 1020 721 1021
rect 722 1020 723 1021
rect 723 1020 724 1021
rect 725 1020 726 1021
rect 720 1021 726 1025
rect 720 1025 721 1026
rect 722 1025 723 1026
rect 723 1025 724 1026
rect 725 1025 726 1026
rect 660 1020 661 1021
rect 662 1020 663 1021
rect 663 1020 664 1021
rect 665 1020 666 1021
rect 660 1021 666 1025
rect 660 1025 661 1026
rect 662 1025 663 1026
rect 663 1025 664 1026
rect 665 1025 666 1026
rect 420 760 421 761
rect 422 760 423 761
rect 423 760 424 761
rect 425 760 426 761
rect 420 761 426 765
rect 420 765 421 766
rect 422 765 423 766
rect 423 765 424 766
rect 425 765 426 766
rect 400 800 401 801
rect 402 800 403 801
rect 403 800 404 801
rect 405 800 406 801
rect 400 801 406 805
rect 400 805 401 806
rect 402 805 403 806
rect 403 805 404 806
rect 405 805 406 806
rect 500 480 501 481
rect 502 480 503 481
rect 503 480 504 481
rect 505 480 506 481
rect 500 481 506 485
rect 500 485 501 486
rect 502 485 503 486
rect 503 485 504 486
rect 505 485 506 486
rect 580 740 581 741
rect 582 740 583 741
rect 583 740 584 741
rect 585 740 586 741
rect 580 741 586 745
rect 580 745 581 746
rect 582 745 583 746
rect 583 745 584 746
rect 585 745 586 746
rect 720 1000 721 1001
rect 722 1000 723 1001
rect 723 1000 724 1001
rect 725 1000 726 1001
rect 720 1001 726 1005
rect 720 1005 721 1006
rect 722 1005 723 1006
rect 723 1005 724 1006
rect 725 1005 726 1006
rect 660 520 661 521
rect 662 520 663 521
rect 663 520 664 521
rect 665 520 666 521
rect 660 521 666 525
rect 660 525 661 526
rect 662 525 663 526
rect 663 525 664 526
rect 665 525 666 526
rect 800 620 801 621
rect 802 620 803 621
rect 803 620 804 621
rect 805 620 806 621
rect 800 621 806 625
rect 800 625 801 626
rect 802 625 803 626
rect 803 625 804 626
rect 805 625 806 626
rect 720 760 721 761
rect 722 760 723 761
rect 723 760 724 761
rect 725 760 726 761
rect 720 761 726 765
rect 720 765 721 766
rect 722 765 723 766
rect 723 765 724 766
rect 725 765 726 766
rect 700 500 701 501
rect 702 500 703 501
rect 703 500 704 501
rect 705 500 706 501
rect 700 501 706 505
rect 700 505 701 506
rect 702 505 703 506
rect 703 505 704 506
rect 705 505 706 506
rect 520 980 521 981
rect 522 980 523 981
rect 523 980 524 981
rect 525 980 526 981
rect 520 981 526 985
rect 520 985 521 986
rect 522 985 523 986
rect 523 985 524 986
rect 525 985 526 986
rect 620 660 621 661
rect 622 660 623 661
rect 623 660 624 661
rect 625 660 626 661
rect 620 661 626 665
rect 620 665 621 666
rect 622 665 623 666
rect 623 665 624 666
rect 625 665 626 666
rect 340 540 341 541
rect 342 540 343 541
rect 343 540 344 541
rect 345 540 346 541
rect 340 541 346 545
rect 340 545 341 546
rect 342 545 343 546
rect 343 545 344 546
rect 345 545 346 546
rect 600 500 601 501
rect 602 500 603 501
rect 603 500 604 501
rect 605 500 606 501
rect 600 501 606 505
rect 600 505 601 506
rect 602 505 603 506
rect 603 505 604 506
rect 605 505 606 506
rect 940 720 941 721
rect 942 720 943 721
rect 943 720 944 721
rect 945 720 946 721
rect 940 721 946 725
rect 940 725 941 726
rect 942 725 943 726
rect 943 725 944 726
rect 945 725 946 726
rect 700 840 701 841
rect 702 840 703 841
rect 703 840 704 841
rect 705 840 706 841
rect 700 841 706 845
rect 700 845 701 846
rect 702 845 703 846
rect 703 845 704 846
rect 705 845 706 846
rect 920 660 921 661
rect 922 660 923 661
rect 923 660 924 661
rect 925 660 926 661
rect 920 661 926 665
rect 920 665 921 666
rect 922 665 923 666
rect 923 665 924 666
rect 925 665 926 666
rect 840 520 841 521
rect 842 520 843 521
rect 843 520 844 521
rect 845 520 846 521
rect 840 521 846 525
rect 840 525 841 526
rect 842 525 843 526
rect 843 525 844 526
rect 845 525 846 526
rect 820 760 821 761
rect 822 760 823 761
rect 823 760 824 761
rect 825 760 826 761
rect 820 761 826 765
rect 820 765 821 766
rect 822 765 823 766
rect 823 765 824 766
rect 825 765 826 766
rect 880 820 881 821
rect 882 820 883 821
rect 883 820 884 821
rect 885 820 886 821
rect 880 821 886 825
rect 880 825 881 826
rect 882 825 883 826
rect 883 825 884 826
rect 885 825 886 826
rect 460 780 461 781
rect 462 780 463 781
rect 463 780 464 781
rect 465 780 466 781
rect 460 781 466 785
rect 460 785 461 786
rect 462 785 463 786
rect 463 785 464 786
rect 465 785 466 786
rect 440 440 441 441
rect 442 440 443 441
rect 443 440 444 441
rect 445 440 446 441
rect 440 441 446 445
rect 440 445 441 446
rect 442 445 443 446
rect 443 445 444 446
rect 445 445 446 446
rect 520 620 521 621
rect 522 620 523 621
rect 523 620 524 621
rect 525 620 526 621
rect 520 621 526 625
rect 520 625 521 626
rect 522 625 523 626
rect 523 625 524 626
rect 525 625 526 626
rect 440 500 441 501
rect 442 500 443 501
rect 443 500 444 501
rect 445 500 446 501
rect 440 501 446 505
rect 440 505 441 506
rect 442 505 443 506
rect 443 505 444 506
rect 445 505 446 506
rect 900 800 901 801
rect 902 800 903 801
rect 903 800 904 801
rect 905 800 906 801
rect 900 801 906 805
rect 900 805 901 806
rect 902 805 903 806
rect 903 805 904 806
rect 905 805 906 806
rect 760 460 761 461
rect 762 460 763 461
rect 763 460 764 461
rect 765 460 766 461
rect 760 461 766 465
rect 760 465 761 466
rect 762 465 763 466
rect 763 465 764 466
rect 765 465 766 466
rect 960 820 961 821
rect 962 820 963 821
rect 963 820 964 821
rect 965 820 966 821
rect 960 821 966 825
rect 960 825 961 826
rect 962 825 963 826
rect 963 825 964 826
rect 965 825 966 826
rect 460 760 461 761
rect 462 760 463 761
rect 463 760 464 761
rect 465 760 466 761
rect 460 761 466 765
rect 460 765 461 766
rect 462 765 463 766
rect 463 765 464 766
rect 465 765 466 766
rect 920 620 921 621
rect 922 620 923 621
rect 923 620 924 621
rect 925 620 926 621
rect 920 621 926 625
rect 920 625 921 626
rect 922 625 923 626
rect 923 625 924 626
rect 925 625 926 626
rect 480 920 481 921
rect 482 920 483 921
rect 483 920 484 921
rect 485 920 486 921
rect 480 921 486 925
rect 480 925 481 926
rect 482 925 483 926
rect 483 925 484 926
rect 485 925 486 926
rect 640 940 641 941
rect 642 940 643 941
rect 643 940 644 941
rect 645 940 646 941
rect 640 941 646 945
rect 640 945 641 946
rect 642 945 643 946
rect 643 945 644 946
rect 645 945 646 946
rect 880 700 881 701
rect 882 700 883 701
rect 883 700 884 701
rect 885 700 886 701
rect 880 701 886 705
rect 880 705 881 706
rect 882 705 883 706
rect 883 705 884 706
rect 885 705 886 706
rect 600 760 601 761
rect 602 760 603 761
rect 603 760 604 761
rect 605 760 606 761
rect 600 761 606 765
rect 600 765 601 766
rect 602 765 603 766
rect 603 765 604 766
rect 605 765 606 766
rect 360 700 361 701
rect 362 700 363 701
rect 363 700 364 701
rect 365 700 366 701
rect 360 701 366 705
rect 360 705 361 706
rect 362 705 363 706
rect 363 705 364 706
rect 365 705 366 706
rect 780 500 781 501
rect 782 500 783 501
rect 783 500 784 501
rect 785 500 786 501
rect 780 501 786 505
rect 780 505 781 506
rect 782 505 783 506
rect 783 505 784 506
rect 785 505 786 506
rect 280 660 281 661
rect 282 660 283 661
rect 283 660 284 661
rect 285 660 286 661
rect 280 661 286 665
rect 280 665 281 666
rect 282 665 283 666
rect 283 665 284 666
rect 285 665 286 666
rect 360 740 361 741
rect 362 740 363 741
rect 363 740 364 741
rect 365 740 366 741
rect 360 741 366 745
rect 360 745 361 746
rect 362 745 363 746
rect 363 745 364 746
rect 365 745 366 746
rect 520 780 521 781
rect 522 780 523 781
rect 523 780 524 781
rect 525 780 526 781
rect 520 781 526 785
rect 520 785 521 786
rect 522 785 523 786
rect 523 785 524 786
rect 525 785 526 786
rect 400 480 401 481
rect 402 480 403 481
rect 403 480 404 481
rect 405 480 406 481
rect 400 481 406 485
rect 400 485 401 486
rect 402 485 403 486
rect 403 485 404 486
rect 405 485 406 486
rect 540 780 541 781
rect 542 780 543 781
rect 543 780 544 781
rect 545 780 546 781
rect 540 781 546 785
rect 540 785 541 786
rect 542 785 543 786
rect 543 785 544 786
rect 545 785 546 786
rect 400 740 401 741
rect 402 740 403 741
rect 403 740 404 741
rect 405 740 406 741
rect 400 741 406 745
rect 400 745 401 746
rect 402 745 403 746
rect 403 745 404 746
rect 405 745 406 746
rect 560 940 561 941
rect 562 940 563 941
rect 563 940 564 941
rect 565 940 566 941
rect 560 941 566 945
rect 560 945 561 946
rect 562 945 563 946
rect 563 945 564 946
rect 565 945 566 946
rect 860 820 861 821
rect 862 820 863 821
rect 863 820 864 821
rect 865 820 866 821
rect 860 821 866 825
rect 860 825 861 826
rect 862 825 863 826
rect 863 825 864 826
rect 865 825 866 826
rect 680 620 681 621
rect 682 620 683 621
rect 683 620 684 621
rect 685 620 686 621
rect 680 621 686 625
rect 680 625 681 626
rect 682 625 683 626
rect 683 625 684 626
rect 685 625 686 626
rect 900 720 901 721
rect 902 720 903 721
rect 903 720 904 721
rect 905 720 906 721
rect 900 721 906 725
rect 900 725 901 726
rect 902 725 903 726
rect 903 725 904 726
rect 905 725 906 726
rect 780 920 781 921
rect 782 920 783 921
rect 783 920 784 921
rect 785 920 786 921
rect 780 921 786 925
rect 780 925 781 926
rect 782 925 783 926
rect 783 925 784 926
rect 785 925 786 926
rect 740 940 741 941
rect 742 940 743 941
rect 743 940 744 941
rect 745 940 746 941
rect 740 941 746 945
rect 740 945 741 946
rect 742 945 743 946
rect 743 945 744 946
rect 745 945 746 946
rect 1000 660 1001 661
rect 1002 660 1003 661
rect 1003 660 1004 661
rect 1005 660 1006 661
rect 1000 661 1006 665
rect 1000 665 1001 666
rect 1002 665 1003 666
rect 1003 665 1004 666
rect 1005 665 1006 666
rect 760 340 761 341
rect 762 340 763 341
rect 763 340 764 341
rect 765 340 766 341
rect 760 341 766 345
rect 760 345 761 346
rect 762 345 763 346
rect 763 345 764 346
rect 765 345 766 346
rect 680 320 681 321
rect 682 320 683 321
rect 683 320 684 321
rect 685 320 686 321
rect 680 321 686 325
rect 680 325 681 326
rect 682 325 683 326
rect 683 325 684 326
rect 685 325 686 326
rect 620 540 621 541
rect 622 540 623 541
rect 623 540 624 541
rect 625 540 626 541
rect 620 541 626 545
rect 620 545 621 546
rect 622 545 623 546
rect 623 545 624 546
rect 625 545 626 546
rect 500 560 501 561
rect 502 560 503 561
rect 503 560 504 561
rect 505 560 506 561
rect 500 561 506 565
rect 500 565 501 566
rect 502 565 503 566
rect 503 565 504 566
rect 505 565 506 566
rect 960 740 961 741
rect 962 740 963 741
rect 963 740 964 741
rect 965 740 966 741
rect 960 741 966 745
rect 960 745 961 746
rect 962 745 963 746
rect 963 745 964 746
rect 965 745 966 746
rect 380 840 381 841
rect 382 840 383 841
rect 383 840 384 841
rect 385 840 386 841
rect 380 841 386 845
rect 380 845 381 846
rect 382 845 383 846
rect 383 845 384 846
rect 385 845 386 846
rect 660 580 661 581
rect 662 580 663 581
rect 663 580 664 581
rect 665 580 666 581
rect 660 581 666 585
rect 660 585 661 586
rect 662 585 663 586
rect 663 585 664 586
rect 665 585 666 586
rect 620 740 621 741
rect 622 740 623 741
rect 623 740 624 741
rect 625 740 626 741
rect 620 741 626 745
rect 620 745 621 746
rect 622 745 623 746
rect 623 745 624 746
rect 625 745 626 746
rect 700 660 701 661
rect 702 660 703 661
rect 703 660 704 661
rect 705 660 706 661
rect 700 661 706 665
rect 700 665 701 666
rect 702 665 703 666
rect 703 665 704 666
rect 705 665 706 666
rect 320 660 321 661
rect 322 660 323 661
rect 323 660 324 661
rect 325 660 326 661
rect 320 661 326 665
rect 320 665 321 666
rect 322 665 323 666
rect 323 665 324 666
rect 325 665 326 666
rect 320 720 321 721
rect 322 720 323 721
rect 323 720 324 721
rect 325 720 326 721
rect 320 721 326 725
rect 320 725 321 726
rect 322 725 323 726
rect 323 725 324 726
rect 325 725 326 726
rect 1040 680 1041 681
rect 1042 680 1043 681
rect 1043 680 1044 681
rect 1045 680 1046 681
rect 1040 681 1046 685
rect 1040 685 1041 686
rect 1042 685 1043 686
rect 1043 685 1044 686
rect 1045 685 1046 686
rect 540 900 541 901
rect 542 900 543 901
rect 543 900 544 901
rect 545 900 546 901
rect 540 901 546 905
rect 540 905 541 906
rect 542 905 543 906
rect 543 905 544 906
rect 545 905 546 906
rect 880 520 881 521
rect 882 520 883 521
rect 883 520 884 521
rect 885 520 886 521
rect 880 521 886 525
rect 880 525 881 526
rect 882 525 883 526
rect 883 525 884 526
rect 885 525 886 526
rect 300 640 301 641
rect 302 640 303 641
rect 303 640 304 641
rect 305 640 306 641
rect 300 641 306 645
rect 300 645 301 646
rect 302 645 303 646
rect 303 645 304 646
rect 305 645 306 646
rect 420 780 421 781
rect 422 780 423 781
rect 423 780 424 781
rect 425 780 426 781
rect 420 781 426 785
rect 420 785 421 786
rect 422 785 423 786
rect 423 785 424 786
rect 425 785 426 786
rect 640 860 641 861
rect 642 860 643 861
rect 643 860 644 861
rect 645 860 646 861
rect 640 861 646 865
rect 640 865 641 866
rect 642 865 643 866
rect 643 865 644 866
rect 645 865 646 866
rect 880 500 881 501
rect 882 500 883 501
rect 883 500 884 501
rect 885 500 886 501
rect 880 501 886 505
rect 880 505 881 506
rect 882 505 883 506
rect 883 505 884 506
rect 885 505 886 506
rect 400 820 401 821
rect 402 820 403 821
rect 403 820 404 821
rect 405 820 406 821
rect 400 821 406 825
rect 400 825 401 826
rect 402 825 403 826
rect 403 825 404 826
rect 405 825 406 826
rect 840 820 841 821
rect 842 820 843 821
rect 843 820 844 821
rect 845 820 846 821
rect 840 821 846 825
rect 840 825 841 826
rect 842 825 843 826
rect 843 825 844 826
rect 845 825 846 826
rect 540 400 541 401
rect 542 400 543 401
rect 543 400 544 401
rect 545 400 546 401
rect 540 401 546 405
rect 540 405 541 406
rect 542 405 543 406
rect 543 405 544 406
rect 545 405 546 406
rect 540 420 541 421
rect 542 420 543 421
rect 543 420 544 421
rect 545 420 546 421
rect 540 421 546 425
rect 540 425 541 426
rect 542 425 543 426
rect 543 425 544 426
rect 545 425 546 426
rect 840 540 841 541
rect 842 540 843 541
rect 843 540 844 541
rect 845 540 846 541
rect 840 541 846 545
rect 840 545 841 546
rect 842 545 843 546
rect 843 545 844 546
rect 845 545 846 546
rect 980 800 981 801
rect 982 800 983 801
rect 983 800 984 801
rect 985 800 986 801
rect 980 801 986 805
rect 980 805 981 806
rect 982 805 983 806
rect 983 805 984 806
rect 985 805 986 806
rect 520 400 521 401
rect 522 400 523 401
rect 523 400 524 401
rect 525 400 526 401
rect 520 401 526 405
rect 520 405 521 406
rect 522 405 523 406
rect 523 405 524 406
rect 525 405 526 406
rect 860 660 861 661
rect 862 660 863 661
rect 863 660 864 661
rect 865 660 866 661
rect 860 661 866 665
rect 860 665 861 666
rect 862 665 863 666
rect 863 665 864 666
rect 865 665 866 666
rect 580 320 581 321
rect 582 320 583 321
rect 583 320 584 321
rect 585 320 586 321
rect 580 321 586 325
rect 580 325 581 326
rect 582 325 583 326
rect 583 325 584 326
rect 585 325 586 326
rect 760 560 761 561
rect 762 560 763 561
rect 763 560 764 561
rect 765 560 766 561
rect 760 561 766 565
rect 760 565 761 566
rect 762 565 763 566
rect 763 565 764 566
rect 765 565 766 566
rect 900 780 901 781
rect 902 780 903 781
rect 903 780 904 781
rect 905 780 906 781
rect 900 781 906 785
rect 900 785 901 786
rect 902 785 903 786
rect 903 785 904 786
rect 905 785 906 786
rect 980 620 981 621
rect 982 620 983 621
rect 983 620 984 621
rect 985 620 986 621
rect 980 621 986 625
rect 980 625 981 626
rect 982 625 983 626
rect 983 625 984 626
rect 985 625 986 626
rect 680 560 681 561
rect 682 560 683 561
rect 683 560 684 561
rect 685 560 686 561
rect 680 561 686 565
rect 680 565 681 566
rect 682 565 683 566
rect 683 565 684 566
rect 685 565 686 566
rect 880 460 881 461
rect 882 460 883 461
rect 883 460 884 461
rect 885 460 886 461
rect 880 461 886 465
rect 880 465 881 466
rect 882 465 883 466
rect 883 465 884 466
rect 885 465 886 466
rect 760 840 761 841
rect 762 840 763 841
rect 763 840 764 841
rect 765 840 766 841
rect 760 841 766 845
rect 760 845 761 846
rect 762 845 763 846
rect 763 845 764 846
rect 765 845 766 846
rect 920 600 921 601
rect 922 600 923 601
rect 923 600 924 601
rect 925 600 926 601
rect 920 601 926 605
rect 920 605 921 606
rect 922 605 923 606
rect 923 605 924 606
rect 925 605 926 606
rect 880 620 881 621
rect 882 620 883 621
rect 883 620 884 621
rect 885 620 886 621
rect 880 621 886 625
rect 880 625 881 626
rect 882 625 883 626
rect 883 625 884 626
rect 885 625 886 626
rect 300 740 301 741
rect 302 740 303 741
rect 303 740 304 741
rect 305 740 306 741
rect 300 741 306 745
rect 300 745 301 746
rect 302 745 303 746
rect 303 745 304 746
rect 305 745 306 746
rect 1020 660 1021 661
rect 1022 660 1023 661
rect 1023 660 1024 661
rect 1025 660 1026 661
rect 1020 661 1026 665
rect 1020 665 1021 666
rect 1022 665 1023 666
rect 1023 665 1024 666
rect 1025 665 1026 666
rect 660 980 661 981
rect 662 980 663 981
rect 663 980 664 981
rect 665 980 666 981
rect 660 981 666 985
rect 660 985 661 986
rect 662 985 663 986
rect 663 985 664 986
rect 665 985 666 986
rect 800 420 801 421
rect 802 420 803 421
rect 803 420 804 421
rect 805 420 806 421
rect 800 421 806 425
rect 800 425 801 426
rect 802 425 803 426
rect 803 425 804 426
rect 805 425 806 426
rect 1000 600 1001 601
rect 1002 600 1003 601
rect 1003 600 1004 601
rect 1005 600 1006 601
rect 1000 601 1006 605
rect 1000 605 1001 606
rect 1002 605 1003 606
rect 1003 605 1004 606
rect 1005 605 1006 606
rect 860 560 861 561
rect 862 560 863 561
rect 863 560 864 561
rect 865 560 866 561
rect 860 561 866 565
rect 860 565 861 566
rect 862 565 863 566
rect 863 565 864 566
rect 865 565 866 566
rect 380 700 381 701
rect 382 700 383 701
rect 383 700 384 701
rect 385 700 386 701
rect 380 701 386 705
rect 380 705 381 706
rect 382 705 383 706
rect 383 705 384 706
rect 385 705 386 706
rect 660 660 661 661
rect 662 660 663 661
rect 663 660 664 661
rect 665 660 666 661
rect 660 661 666 665
rect 660 665 661 666
rect 662 665 663 666
rect 663 665 664 666
rect 665 665 666 666
rect 520 940 521 941
rect 522 940 523 941
rect 523 940 524 941
rect 525 940 526 941
rect 520 941 526 945
rect 520 945 521 946
rect 522 945 523 946
rect 523 945 524 946
rect 525 945 526 946
rect 740 800 741 801
rect 742 800 743 801
rect 743 800 744 801
rect 745 800 746 801
rect 740 801 746 805
rect 740 805 741 806
rect 742 805 743 806
rect 743 805 744 806
rect 745 805 746 806
rect 520 500 521 501
rect 522 500 523 501
rect 523 500 524 501
rect 525 500 526 501
rect 520 501 526 505
rect 520 505 521 506
rect 522 505 523 506
rect 523 505 524 506
rect 525 505 526 506
rect 540 480 541 481
rect 542 480 543 481
rect 543 480 544 481
rect 545 480 546 481
rect 540 481 546 485
rect 540 485 541 486
rect 542 485 543 486
rect 543 485 544 486
rect 545 485 546 486
rect 400 580 401 581
rect 402 580 403 581
rect 403 580 404 581
rect 405 580 406 581
rect 400 581 406 585
rect 400 585 401 586
rect 402 585 403 586
rect 403 585 404 586
rect 405 585 406 586
rect 980 640 981 641
rect 982 640 983 641
rect 983 640 984 641
rect 985 640 986 641
rect 980 641 986 645
rect 980 645 981 646
rect 982 645 983 646
rect 983 645 984 646
rect 985 645 986 646
rect 460 820 461 821
rect 462 820 463 821
rect 463 820 464 821
rect 465 820 466 821
rect 460 821 466 825
rect 460 825 461 826
rect 462 825 463 826
rect 463 825 464 826
rect 465 825 466 826
rect 580 480 581 481
rect 582 480 583 481
rect 583 480 584 481
rect 585 480 586 481
rect 580 481 586 485
rect 580 485 581 486
rect 582 485 583 486
rect 583 485 584 486
rect 585 485 586 486
rect 420 580 421 581
rect 422 580 423 581
rect 423 580 424 581
rect 425 580 426 581
rect 420 581 426 585
rect 420 585 421 586
rect 422 585 423 586
rect 423 585 424 586
rect 425 585 426 586
rect 400 780 401 781
rect 402 780 403 781
rect 403 780 404 781
rect 405 780 406 781
rect 400 781 406 785
rect 400 785 401 786
rect 402 785 403 786
rect 403 785 404 786
rect 405 785 406 786
rect 300 800 301 801
rect 302 800 303 801
rect 303 800 304 801
rect 305 800 306 801
rect 300 801 306 805
rect 300 805 301 806
rect 302 805 303 806
rect 303 805 304 806
rect 305 805 306 806
rect 940 520 941 521
rect 942 520 943 521
rect 943 520 944 521
rect 945 520 946 521
rect 940 521 946 525
rect 940 525 941 526
rect 942 525 943 526
rect 943 525 944 526
rect 945 525 946 526
rect 580 1000 581 1001
rect 582 1000 583 1001
rect 583 1000 584 1001
rect 585 1000 586 1001
rect 580 1001 586 1005
rect 580 1005 581 1006
rect 582 1005 583 1006
rect 583 1005 584 1006
rect 585 1005 586 1006
rect 680 280 681 281
rect 682 280 683 281
rect 683 280 684 281
rect 685 280 686 281
rect 680 281 686 285
rect 680 285 681 286
rect 682 285 683 286
rect 683 285 684 286
rect 685 285 686 286
rect 880 440 881 441
rect 882 440 883 441
rect 883 440 884 441
rect 885 440 886 441
rect 880 441 886 445
rect 880 445 881 446
rect 882 445 883 446
rect 883 445 884 446
rect 885 445 886 446
rect 400 600 401 601
rect 402 600 403 601
rect 403 600 404 601
rect 405 600 406 601
rect 400 601 406 605
rect 400 605 401 606
rect 402 605 403 606
rect 403 605 404 606
rect 405 605 406 606
rect 900 560 901 561
rect 902 560 903 561
rect 903 560 904 561
rect 905 560 906 561
rect 900 561 906 565
rect 900 565 901 566
rect 902 565 903 566
rect 903 565 904 566
rect 905 565 906 566
rect 1000 760 1001 761
rect 1002 760 1003 761
rect 1003 760 1004 761
rect 1005 760 1006 761
rect 1000 761 1006 765
rect 1000 765 1001 766
rect 1002 765 1003 766
rect 1003 765 1004 766
rect 1005 765 1006 766
rect 320 640 321 641
rect 322 640 323 641
rect 323 640 324 641
rect 325 640 326 641
rect 320 641 326 645
rect 320 645 321 646
rect 322 645 323 646
rect 323 645 324 646
rect 325 645 326 646
rect 680 880 681 881
rect 682 880 683 881
rect 683 880 684 881
rect 685 880 686 881
rect 680 881 686 885
rect 680 885 681 886
rect 682 885 683 886
rect 683 885 684 886
rect 685 885 686 886
rect 860 800 861 801
rect 862 800 863 801
rect 863 800 864 801
rect 865 800 866 801
rect 860 801 866 805
rect 860 805 861 806
rect 862 805 863 806
rect 863 805 864 806
rect 865 805 866 806
rect 860 700 861 701
rect 862 700 863 701
rect 863 700 864 701
rect 865 700 866 701
rect 860 701 866 705
rect 860 705 861 706
rect 862 705 863 706
rect 863 705 864 706
rect 865 705 866 706
rect 1000 680 1001 681
rect 1002 680 1003 681
rect 1003 680 1004 681
rect 1005 680 1006 681
rect 1000 681 1006 685
rect 1000 685 1001 686
rect 1002 685 1003 686
rect 1003 685 1004 686
rect 1005 685 1006 686
rect 740 700 741 701
rect 742 700 743 701
rect 743 700 744 701
rect 745 700 746 701
rect 740 701 746 705
rect 740 705 741 706
rect 742 705 743 706
rect 743 705 744 706
rect 745 705 746 706
rect 300 680 301 681
rect 302 680 303 681
rect 303 680 304 681
rect 305 680 306 681
rect 300 681 306 685
rect 300 685 301 686
rect 302 685 303 686
rect 303 685 304 686
rect 305 685 306 686
rect 680 760 681 761
rect 682 760 683 761
rect 683 760 684 761
rect 685 760 686 761
rect 680 761 686 765
rect 680 765 681 766
rect 682 765 683 766
rect 683 765 684 766
rect 685 765 686 766
rect 660 400 661 401
rect 662 400 663 401
rect 663 400 664 401
rect 665 400 666 401
rect 660 401 666 405
rect 660 405 661 406
rect 662 405 663 406
rect 663 405 664 406
rect 665 405 666 406
rect 380 720 381 721
rect 382 720 383 721
rect 383 720 384 721
rect 385 720 386 721
rect 380 721 386 725
rect 380 725 381 726
rect 382 725 383 726
rect 383 725 384 726
rect 385 725 386 726
rect 300 720 301 721
rect 302 720 303 721
rect 303 720 304 721
rect 305 720 306 721
rect 300 721 306 725
rect 300 725 301 726
rect 302 725 303 726
rect 303 725 304 726
rect 305 725 306 726
rect 700 980 701 981
rect 702 980 703 981
rect 703 980 704 981
rect 705 980 706 981
rect 700 981 706 985
rect 700 985 701 986
rect 702 985 703 986
rect 703 985 704 986
rect 705 985 706 986
rect 540 740 541 741
rect 542 740 543 741
rect 543 740 544 741
rect 545 740 546 741
rect 540 741 546 745
rect 540 745 541 746
rect 542 745 543 746
rect 543 745 544 746
rect 545 745 546 746
rect 820 720 821 721
rect 822 720 823 721
rect 823 720 824 721
rect 825 720 826 721
rect 820 721 826 725
rect 820 725 821 726
rect 822 725 823 726
rect 823 725 824 726
rect 825 725 826 726
rect 640 760 641 761
rect 642 760 643 761
rect 643 760 644 761
rect 645 760 646 761
rect 640 761 646 765
rect 640 765 641 766
rect 642 765 643 766
rect 643 765 644 766
rect 645 765 646 766
rect 760 600 761 601
rect 762 600 763 601
rect 763 600 764 601
rect 765 600 766 601
rect 760 601 766 605
rect 760 605 761 606
rect 762 605 763 606
rect 763 605 764 606
rect 765 605 766 606
rect 840 580 841 581
rect 842 580 843 581
rect 843 580 844 581
rect 845 580 846 581
rect 840 581 846 585
rect 840 585 841 586
rect 842 585 843 586
rect 843 585 844 586
rect 845 585 846 586
rect 420 600 421 601
rect 422 600 423 601
rect 423 600 424 601
rect 425 600 426 601
rect 420 601 426 605
rect 420 605 421 606
rect 422 605 423 606
rect 423 605 424 606
rect 425 605 426 606
rect 740 440 741 441
rect 742 440 743 441
rect 743 440 744 441
rect 745 440 746 441
rect 740 441 746 445
rect 740 445 741 446
rect 742 445 743 446
rect 743 445 744 446
rect 745 445 746 446
rect 800 960 801 961
rect 802 960 803 961
rect 803 960 804 961
rect 805 960 806 961
rect 800 961 806 965
rect 800 965 801 966
rect 802 965 803 966
rect 803 965 804 966
rect 805 965 806 966
rect 780 860 781 861
rect 782 860 783 861
rect 783 860 784 861
rect 785 860 786 861
rect 780 861 786 865
rect 780 865 781 866
rect 782 865 783 866
rect 783 865 784 866
rect 785 865 786 866
rect 680 1020 681 1021
rect 682 1020 683 1021
rect 683 1020 684 1021
rect 685 1020 686 1021
rect 680 1021 686 1025
rect 680 1025 681 1026
rect 682 1025 683 1026
rect 683 1025 684 1026
rect 685 1025 686 1026
rect 540 960 541 961
rect 542 960 543 961
rect 543 960 544 961
rect 545 960 546 961
rect 540 961 546 965
rect 540 965 541 966
rect 542 965 543 966
rect 543 965 544 966
rect 545 965 546 966
rect 980 600 981 601
rect 982 600 983 601
rect 983 600 984 601
rect 985 600 986 601
rect 980 601 986 605
rect 980 605 981 606
rect 982 605 983 606
rect 983 605 984 606
rect 985 605 986 606
rect 800 920 801 921
rect 802 920 803 921
rect 803 920 804 921
rect 805 920 806 921
rect 800 921 806 925
rect 800 925 801 926
rect 802 925 803 926
rect 803 925 804 926
rect 805 925 806 926
rect 960 660 961 661
rect 962 660 963 661
rect 963 660 964 661
rect 965 660 966 661
rect 960 661 966 665
rect 960 665 961 666
rect 962 665 963 666
rect 963 665 964 666
rect 965 665 966 666
rect 640 1000 641 1001
rect 642 1000 643 1001
rect 643 1000 644 1001
rect 645 1000 646 1001
rect 640 1001 646 1005
rect 640 1005 641 1006
rect 642 1005 643 1006
rect 643 1005 644 1006
rect 645 1005 646 1006
rect 320 580 321 581
rect 322 580 323 581
rect 323 580 324 581
rect 325 580 326 581
rect 320 581 326 585
rect 320 585 321 586
rect 322 585 323 586
rect 323 585 324 586
rect 325 585 326 586
rect 580 340 581 341
rect 582 340 583 341
rect 583 340 584 341
rect 585 340 586 341
rect 580 341 586 345
rect 580 345 581 346
rect 582 345 583 346
rect 583 345 584 346
rect 585 345 586 346
rect 580 820 581 821
rect 582 820 583 821
rect 583 820 584 821
rect 585 820 586 821
rect 580 821 586 825
rect 580 825 581 826
rect 582 825 583 826
rect 583 825 584 826
rect 585 825 586 826
rect 760 820 761 821
rect 762 820 763 821
rect 763 820 764 821
rect 765 820 766 821
rect 760 821 766 825
rect 760 825 761 826
rect 762 825 763 826
rect 763 825 764 826
rect 765 825 766 826
rect 580 860 581 861
rect 582 860 583 861
rect 583 860 584 861
rect 585 860 586 861
rect 580 861 586 865
rect 580 865 581 866
rect 582 865 583 866
rect 583 865 584 866
rect 585 865 586 866
rect 700 620 701 621
rect 702 620 703 621
rect 703 620 704 621
rect 705 620 706 621
rect 700 621 706 625
rect 700 625 701 626
rect 702 625 703 626
rect 703 625 704 626
rect 705 625 706 626
rect 520 600 521 601
rect 522 600 523 601
rect 523 600 524 601
rect 525 600 526 601
rect 520 601 526 605
rect 520 605 521 606
rect 522 605 523 606
rect 523 605 524 606
rect 525 605 526 606
rect 580 920 581 921
rect 582 920 583 921
rect 583 920 584 921
rect 585 920 586 921
rect 580 921 586 925
rect 580 925 581 926
rect 582 925 583 926
rect 583 925 584 926
rect 585 925 586 926
rect 880 660 881 661
rect 882 660 883 661
rect 883 660 884 661
rect 885 660 886 661
rect 880 661 886 665
rect 880 665 881 666
rect 882 665 883 666
rect 883 665 884 666
rect 885 665 886 666
rect 460 880 461 881
rect 462 880 463 881
rect 463 880 464 881
rect 465 880 466 881
rect 460 881 466 885
rect 460 885 461 886
rect 462 885 463 886
rect 463 885 464 886
rect 465 885 466 886
rect 520 900 521 901
rect 522 900 523 901
rect 523 900 524 901
rect 525 900 526 901
rect 520 901 526 905
rect 520 905 521 906
rect 522 905 523 906
rect 523 905 524 906
rect 525 905 526 906
rect 880 680 881 681
rect 882 680 883 681
rect 883 680 884 681
rect 885 680 886 681
rect 880 681 886 685
rect 880 685 881 686
rect 882 685 883 686
rect 883 685 884 686
rect 885 685 886 686
rect 440 780 441 781
rect 442 780 443 781
rect 443 780 444 781
rect 445 780 446 781
rect 440 781 446 785
rect 440 785 441 786
rect 442 785 443 786
rect 443 785 444 786
rect 445 785 446 786
rect 400 860 401 861
rect 402 860 403 861
rect 403 860 404 861
rect 405 860 406 861
rect 400 861 406 865
rect 400 865 401 866
rect 402 865 403 866
rect 403 865 404 866
rect 405 865 406 866
rect 680 960 681 961
rect 682 960 683 961
rect 683 960 684 961
rect 685 960 686 961
rect 680 961 686 965
rect 680 965 681 966
rect 682 965 683 966
rect 683 965 684 966
rect 685 965 686 966
rect 820 460 821 461
rect 822 460 823 461
rect 823 460 824 461
rect 825 460 826 461
rect 820 461 826 465
rect 820 465 821 466
rect 822 465 823 466
rect 823 465 824 466
rect 825 465 826 466
rect 720 500 721 501
rect 722 500 723 501
rect 723 500 724 501
rect 725 500 726 501
rect 720 501 726 505
rect 720 505 721 506
rect 722 505 723 506
rect 723 505 724 506
rect 725 505 726 506
rect 500 820 501 821
rect 502 820 503 821
rect 503 820 504 821
rect 505 820 506 821
rect 500 821 506 825
rect 500 825 501 826
rect 502 825 503 826
rect 503 825 504 826
rect 505 825 506 826
rect 440 800 441 801
rect 442 800 443 801
rect 443 800 444 801
rect 445 800 446 801
rect 440 801 446 805
rect 440 805 441 806
rect 442 805 443 806
rect 443 805 444 806
rect 445 805 446 806
rect 760 740 761 741
rect 762 740 763 741
rect 763 740 764 741
rect 765 740 766 741
rect 760 741 766 745
rect 760 745 761 746
rect 762 745 763 746
rect 763 745 764 746
rect 765 745 766 746
rect 900 660 901 661
rect 902 660 903 661
rect 903 660 904 661
rect 905 660 906 661
rect 900 661 906 665
rect 900 665 901 666
rect 902 665 903 666
rect 903 665 904 666
rect 905 665 906 666
rect 560 800 561 801
rect 562 800 563 801
rect 563 800 564 801
rect 565 800 566 801
rect 560 801 566 805
rect 560 805 561 806
rect 562 805 563 806
rect 563 805 564 806
rect 565 805 566 806
rect 920 820 921 821
rect 922 820 923 821
rect 923 820 924 821
rect 925 820 926 821
rect 920 821 926 825
rect 920 825 921 826
rect 922 825 923 826
rect 923 825 924 826
rect 925 825 926 826
rect 380 740 381 741
rect 382 740 383 741
rect 383 740 384 741
rect 385 740 386 741
rect 380 741 386 745
rect 380 745 381 746
rect 382 745 383 746
rect 383 745 384 746
rect 385 745 386 746
rect 660 700 661 701
rect 662 700 663 701
rect 663 700 664 701
rect 665 700 666 701
rect 660 701 666 705
rect 660 705 661 706
rect 662 705 663 706
rect 663 705 664 706
rect 665 705 666 706
rect 540 840 541 841
rect 542 840 543 841
rect 543 840 544 841
rect 545 840 546 841
rect 540 841 546 845
rect 540 845 541 846
rect 542 845 543 846
rect 543 845 544 846
rect 545 845 546 846
rect 300 580 301 581
rect 302 580 303 581
rect 303 580 304 581
rect 305 580 306 581
rect 300 581 306 585
rect 300 585 301 586
rect 302 585 303 586
rect 303 585 304 586
rect 305 585 306 586
rect 780 700 781 701
rect 782 700 783 701
rect 783 700 784 701
rect 785 700 786 701
rect 780 701 786 705
rect 780 705 781 706
rect 782 705 783 706
rect 783 705 784 706
rect 785 705 786 706
rect 480 900 481 901
rect 482 900 483 901
rect 483 900 484 901
rect 485 900 486 901
rect 480 901 486 905
rect 480 905 481 906
rect 482 905 483 906
rect 483 905 484 906
rect 485 905 486 906
rect 740 1000 741 1001
rect 742 1000 743 1001
rect 743 1000 744 1001
rect 745 1000 746 1001
rect 740 1001 746 1005
rect 740 1005 741 1006
rect 742 1005 743 1006
rect 743 1005 744 1006
rect 745 1005 746 1006
rect 660 480 661 481
rect 662 480 663 481
rect 663 480 664 481
rect 665 480 666 481
rect 660 481 666 485
rect 660 485 661 486
rect 662 485 663 486
rect 663 485 664 486
rect 665 485 666 486
rect 480 720 481 721
rect 482 720 483 721
rect 483 720 484 721
rect 485 720 486 721
rect 480 721 486 725
rect 480 725 481 726
rect 482 725 483 726
rect 483 725 484 726
rect 485 725 486 726
rect 860 580 861 581
rect 862 580 863 581
rect 863 580 864 581
rect 865 580 866 581
rect 860 581 866 585
rect 860 585 861 586
rect 862 585 863 586
rect 863 585 864 586
rect 865 585 866 586
rect 420 500 421 501
rect 422 500 423 501
rect 423 500 424 501
rect 425 500 426 501
rect 420 501 426 505
rect 420 505 421 506
rect 422 505 423 506
rect 423 505 424 506
rect 425 505 426 506
rect 500 500 501 501
rect 502 500 503 501
rect 503 500 504 501
rect 505 500 506 501
rect 500 501 506 505
rect 500 505 501 506
rect 502 505 503 506
rect 503 505 504 506
rect 505 505 506 506
rect 640 680 641 681
rect 642 680 643 681
rect 643 680 644 681
rect 645 680 646 681
rect 640 681 646 685
rect 640 685 641 686
rect 642 685 643 686
rect 643 685 644 686
rect 645 685 646 686
rect 900 740 901 741
rect 902 740 903 741
rect 903 740 904 741
rect 905 740 906 741
rect 900 741 906 745
rect 900 745 901 746
rect 902 745 903 746
rect 903 745 904 746
rect 905 745 906 746
rect 600 960 601 961
rect 602 960 603 961
rect 603 960 604 961
rect 605 960 606 961
rect 600 961 606 965
rect 600 965 601 966
rect 602 965 603 966
rect 603 965 604 966
rect 605 965 606 966
rect 660 720 661 721
rect 662 720 663 721
rect 663 720 664 721
rect 665 720 666 721
rect 660 721 666 725
rect 660 725 661 726
rect 662 725 663 726
rect 663 725 664 726
rect 665 725 666 726
rect 780 800 781 801
rect 782 800 783 801
rect 783 800 784 801
rect 785 800 786 801
rect 780 801 786 805
rect 780 805 781 806
rect 782 805 783 806
rect 783 805 784 806
rect 785 805 786 806
rect 840 760 841 761
rect 842 760 843 761
rect 843 760 844 761
rect 845 760 846 761
rect 840 761 846 765
rect 840 765 841 766
rect 842 765 843 766
rect 843 765 844 766
rect 845 765 846 766
rect 620 820 621 821
rect 622 820 623 821
rect 623 820 624 821
rect 625 820 626 821
rect 620 821 626 825
rect 620 825 621 826
rect 622 825 623 826
rect 623 825 624 826
rect 625 825 626 826
rect 380 660 381 661
rect 382 660 383 661
rect 383 660 384 661
rect 385 660 386 661
rect 380 661 386 665
rect 380 665 381 666
rect 382 665 383 666
rect 383 665 384 666
rect 385 665 386 666
rect 720 700 721 701
rect 722 700 723 701
rect 723 700 724 701
rect 725 700 726 701
rect 720 701 726 705
rect 720 705 721 706
rect 722 705 723 706
rect 723 705 724 706
rect 725 705 726 706
rect 760 760 761 761
rect 762 760 763 761
rect 763 760 764 761
rect 765 760 766 761
rect 760 761 766 765
rect 760 765 761 766
rect 762 765 763 766
rect 763 765 764 766
rect 765 765 766 766
rect 640 440 641 441
rect 642 440 643 441
rect 643 440 644 441
rect 645 440 646 441
rect 640 441 646 445
rect 640 445 641 446
rect 642 445 643 446
rect 643 445 644 446
rect 645 445 646 446
rect 820 420 821 421
rect 822 420 823 421
rect 823 420 824 421
rect 825 420 826 421
rect 820 421 826 425
rect 820 425 821 426
rect 822 425 823 426
rect 823 425 824 426
rect 825 425 826 426
rect 440 660 441 661
rect 442 660 443 661
rect 443 660 444 661
rect 445 660 446 661
rect 440 661 446 665
rect 440 665 441 666
rect 442 665 443 666
rect 443 665 444 666
rect 445 665 446 666
rect 780 620 781 621
rect 782 620 783 621
rect 783 620 784 621
rect 785 620 786 621
rect 780 621 786 625
rect 780 625 781 626
rect 782 625 783 626
rect 783 625 784 626
rect 785 625 786 626
rect 280 680 281 681
rect 282 680 283 681
rect 283 680 284 681
rect 285 680 286 681
rect 280 681 286 685
rect 280 685 281 686
rect 282 685 283 686
rect 283 685 284 686
rect 285 685 286 686
rect 740 920 741 921
rect 742 920 743 921
rect 743 920 744 921
rect 745 920 746 921
rect 740 921 746 925
rect 740 925 741 926
rect 742 925 743 926
rect 743 925 744 926
rect 745 925 746 926
rect 420 560 421 561
rect 422 560 423 561
rect 423 560 424 561
rect 425 560 426 561
rect 420 561 426 565
rect 420 565 421 566
rect 422 565 423 566
rect 423 565 424 566
rect 425 565 426 566
rect 460 800 461 801
rect 462 800 463 801
rect 463 800 464 801
rect 465 800 466 801
rect 460 801 466 805
rect 460 805 461 806
rect 462 805 463 806
rect 463 805 464 806
rect 465 805 466 806
rect 460 480 461 481
rect 462 480 463 481
rect 463 480 464 481
rect 465 480 466 481
rect 460 481 466 485
rect 460 485 461 486
rect 462 485 463 486
rect 463 485 464 486
rect 465 485 466 486
rect 840 640 841 641
rect 842 640 843 641
rect 843 640 844 641
rect 845 640 846 641
rect 840 641 846 645
rect 840 645 841 646
rect 842 645 843 646
rect 843 645 844 646
rect 845 645 846 646
rect 360 780 361 781
rect 362 780 363 781
rect 363 780 364 781
rect 365 780 366 781
rect 360 781 366 785
rect 360 785 361 786
rect 362 785 363 786
rect 363 785 364 786
rect 365 785 366 786
rect 620 940 621 941
rect 622 940 623 941
rect 623 940 624 941
rect 625 940 626 941
rect 620 941 626 945
rect 620 945 621 946
rect 622 945 623 946
rect 623 945 624 946
rect 625 945 626 946
rect 880 740 881 741
rect 882 740 883 741
rect 883 740 884 741
rect 885 740 886 741
rect 880 741 886 745
rect 880 745 881 746
rect 882 745 883 746
rect 883 745 884 746
rect 885 745 886 746
rect 820 940 821 941
rect 822 940 823 941
rect 823 940 824 941
rect 825 940 826 941
rect 820 941 826 945
rect 820 945 821 946
rect 822 945 823 946
rect 823 945 824 946
rect 825 945 826 946
rect 600 860 601 861
rect 602 860 603 861
rect 603 860 604 861
rect 605 860 606 861
rect 600 861 606 865
rect 600 865 601 866
rect 602 865 603 866
rect 603 865 604 866
rect 605 865 606 866
rect 680 820 681 821
rect 682 820 683 821
rect 683 820 684 821
rect 685 820 686 821
rect 680 821 686 825
rect 680 825 681 826
rect 682 825 683 826
rect 683 825 684 826
rect 685 825 686 826
rect 820 580 821 581
rect 822 580 823 581
rect 823 580 824 581
rect 825 580 826 581
rect 820 581 826 585
rect 820 585 821 586
rect 822 585 823 586
rect 823 585 824 586
rect 825 585 826 586
rect 620 620 621 621
rect 622 620 623 621
rect 623 620 624 621
rect 625 620 626 621
rect 620 621 626 625
rect 620 625 621 626
rect 622 625 623 626
rect 623 625 624 626
rect 625 625 626 626
rect 600 880 601 881
rect 602 880 603 881
rect 603 880 604 881
rect 605 880 606 881
rect 600 881 606 885
rect 600 885 601 886
rect 602 885 603 886
rect 603 885 604 886
rect 605 885 606 886
rect 380 500 381 501
rect 382 500 383 501
rect 383 500 384 501
rect 385 500 386 501
rect 380 501 386 505
rect 380 505 381 506
rect 382 505 383 506
rect 383 505 384 506
rect 385 505 386 506
rect 580 500 581 501
rect 582 500 583 501
rect 583 500 584 501
rect 585 500 586 501
rect 580 501 586 505
rect 580 505 581 506
rect 582 505 583 506
rect 583 505 584 506
rect 585 505 586 506
rect 880 800 881 801
rect 882 800 883 801
rect 883 800 884 801
rect 885 800 886 801
rect 880 801 886 805
rect 880 805 881 806
rect 882 805 883 806
rect 883 805 884 806
rect 885 805 886 806
rect 580 520 581 521
rect 582 520 583 521
rect 583 520 584 521
rect 585 520 586 521
rect 580 521 586 525
rect 580 525 581 526
rect 582 525 583 526
rect 583 525 584 526
rect 585 525 586 526
rect 880 780 881 781
rect 882 780 883 781
rect 883 780 884 781
rect 885 780 886 781
rect 880 781 886 785
rect 880 785 881 786
rect 882 785 883 786
rect 883 785 884 786
rect 885 785 886 786
rect 520 380 521 381
rect 522 380 523 381
rect 523 380 524 381
rect 525 380 526 381
rect 520 381 526 385
rect 520 385 521 386
rect 522 385 523 386
rect 523 385 524 386
rect 525 385 526 386
rect 880 880 881 881
rect 882 880 883 881
rect 883 880 884 881
rect 885 880 886 881
rect 880 881 886 885
rect 880 885 881 886
rect 882 885 883 886
rect 883 885 884 886
rect 885 885 886 886
rect 460 700 461 701
rect 462 700 463 701
rect 463 700 464 701
rect 465 700 466 701
rect 460 701 466 705
rect 460 705 461 706
rect 462 705 463 706
rect 463 705 464 706
rect 465 705 466 706
rect 280 640 281 641
rect 282 640 283 641
rect 283 640 284 641
rect 285 640 286 641
rect 280 641 286 645
rect 280 645 281 646
rect 282 645 283 646
rect 283 645 284 646
rect 285 645 286 646
rect 700 440 701 441
rect 702 440 703 441
rect 703 440 704 441
rect 705 440 706 441
rect 700 441 706 445
rect 700 445 701 446
rect 702 445 703 446
rect 703 445 704 446
rect 705 445 706 446
rect 640 360 641 361
rect 642 360 643 361
rect 643 360 644 361
rect 645 360 646 361
rect 640 361 646 365
rect 640 365 641 366
rect 642 365 643 366
rect 643 365 644 366
rect 645 365 646 366
rect 860 720 861 721
rect 862 720 863 721
rect 863 720 864 721
rect 865 720 866 721
rect 860 721 866 725
rect 860 725 861 726
rect 862 725 863 726
rect 863 725 864 726
rect 865 725 866 726
rect 960 780 961 781
rect 962 780 963 781
rect 963 780 964 781
rect 965 780 966 781
rect 960 781 966 785
rect 960 785 961 786
rect 962 785 963 786
rect 963 785 964 786
rect 965 785 966 786
rect 1020 720 1021 721
rect 1022 720 1023 721
rect 1023 720 1024 721
rect 1025 720 1026 721
rect 1020 721 1026 725
rect 1020 725 1021 726
rect 1022 725 1023 726
rect 1023 725 1024 726
rect 1025 725 1026 726
rect 880 840 881 841
rect 882 840 883 841
rect 883 840 884 841
rect 885 840 886 841
rect 880 841 886 845
rect 880 845 881 846
rect 882 845 883 846
rect 883 845 884 846
rect 885 845 886 846
rect 640 420 641 421
rect 642 420 643 421
rect 643 420 644 421
rect 645 420 646 421
rect 640 421 646 425
rect 640 425 641 426
rect 642 425 643 426
rect 643 425 644 426
rect 645 425 646 426
rect 840 600 841 601
rect 842 600 843 601
rect 843 600 844 601
rect 845 600 846 601
rect 840 601 846 605
rect 840 605 841 606
rect 842 605 843 606
rect 843 605 844 606
rect 845 605 846 606
rect 560 560 561 561
rect 562 560 563 561
rect 563 560 564 561
rect 565 560 566 561
rect 560 561 566 565
rect 560 565 561 566
rect 562 565 563 566
rect 563 565 564 566
rect 565 565 566 566
rect 740 900 741 901
rect 742 900 743 901
rect 743 900 744 901
rect 745 900 746 901
rect 740 901 746 905
rect 740 905 741 906
rect 742 905 743 906
rect 743 905 744 906
rect 745 905 746 906
rect 580 960 581 961
rect 582 960 583 961
rect 583 960 584 961
rect 585 960 586 961
rect 580 961 586 965
rect 580 965 581 966
rect 582 965 583 966
rect 583 965 584 966
rect 585 965 586 966
rect 500 900 501 901
rect 502 900 503 901
rect 503 900 504 901
rect 505 900 506 901
rect 500 901 506 905
rect 500 905 501 906
rect 502 905 503 906
rect 503 905 504 906
rect 505 905 506 906
rect 460 520 461 521
rect 462 520 463 521
rect 463 520 464 521
rect 465 520 466 521
rect 460 521 466 525
rect 460 525 461 526
rect 462 525 463 526
rect 463 525 464 526
rect 465 525 466 526
rect 680 580 681 581
rect 682 580 683 581
rect 683 580 684 581
rect 685 580 686 581
rect 680 581 686 585
rect 680 585 681 586
rect 682 585 683 586
rect 683 585 684 586
rect 685 585 686 586
rect 940 680 941 681
rect 942 680 943 681
rect 943 680 944 681
rect 945 680 946 681
rect 940 681 946 685
rect 940 685 941 686
rect 942 685 943 686
rect 943 685 944 686
rect 945 685 946 686
rect 900 520 901 521
rect 902 520 903 521
rect 903 520 904 521
rect 905 520 906 521
rect 900 521 906 525
rect 900 525 901 526
rect 902 525 903 526
rect 903 525 904 526
rect 905 525 906 526
rect 600 400 601 401
rect 602 400 603 401
rect 603 400 604 401
rect 605 400 606 401
rect 600 401 606 405
rect 600 405 601 406
rect 602 405 603 406
rect 603 405 604 406
rect 605 405 606 406
rect 580 440 581 441
rect 582 440 583 441
rect 583 440 584 441
rect 585 440 586 441
rect 580 441 586 445
rect 580 445 581 446
rect 582 445 583 446
rect 583 445 584 446
rect 585 445 586 446
rect 560 500 561 501
rect 562 500 563 501
rect 563 500 564 501
rect 565 500 566 501
rect 560 501 566 505
rect 560 505 561 506
rect 562 505 563 506
rect 563 505 564 506
rect 565 505 566 506
rect 500 860 501 861
rect 502 860 503 861
rect 503 860 504 861
rect 505 860 506 861
rect 500 861 506 865
rect 500 865 501 866
rect 502 865 503 866
rect 503 865 504 866
rect 505 865 506 866
rect 480 820 481 821
rect 482 820 483 821
rect 483 820 484 821
rect 485 820 486 821
rect 480 821 486 825
rect 480 825 481 826
rect 482 825 483 826
rect 483 825 484 826
rect 485 825 486 826
rect 720 860 721 861
rect 722 860 723 861
rect 723 860 724 861
rect 725 860 726 861
rect 720 861 726 865
rect 720 865 721 866
rect 722 865 723 866
rect 723 865 724 866
rect 725 865 726 866
rect 600 440 601 441
rect 602 440 603 441
rect 603 440 604 441
rect 605 440 606 441
rect 600 441 606 445
rect 600 445 601 446
rect 602 445 603 446
rect 603 445 604 446
rect 605 445 606 446
rect 820 540 821 541
rect 822 540 823 541
rect 823 540 824 541
rect 825 540 826 541
rect 820 541 826 545
rect 820 545 821 546
rect 822 545 823 546
rect 823 545 824 546
rect 825 545 826 546
rect 660 360 661 361
rect 662 360 663 361
rect 663 360 664 361
rect 665 360 666 361
rect 660 361 666 365
rect 660 365 661 366
rect 662 365 663 366
rect 663 365 664 366
rect 665 365 666 366
rect 580 760 581 761
rect 582 760 583 761
rect 583 760 584 761
rect 585 760 586 761
rect 580 761 586 765
rect 580 765 581 766
rect 582 765 583 766
rect 583 765 584 766
rect 585 765 586 766
rect 600 940 601 941
rect 602 940 603 941
rect 603 940 604 941
rect 605 940 606 941
rect 600 941 606 945
rect 600 945 601 946
rect 602 945 603 946
rect 603 945 604 946
rect 605 945 606 946
rect 520 700 521 701
rect 522 700 523 701
rect 523 700 524 701
rect 525 700 526 701
rect 520 701 526 705
rect 520 705 521 706
rect 522 705 523 706
rect 523 705 524 706
rect 525 705 526 706
rect 680 500 681 501
rect 682 500 683 501
rect 683 500 684 501
rect 685 500 686 501
rect 680 501 686 505
rect 680 505 681 506
rect 682 505 683 506
rect 683 505 684 506
rect 685 505 686 506
rect 780 680 781 681
rect 782 680 783 681
rect 783 680 784 681
rect 785 680 786 681
rect 780 681 786 685
rect 780 685 781 686
rect 782 685 783 686
rect 783 685 784 686
rect 785 685 786 686
rect 280 600 281 601
rect 282 600 283 601
rect 283 600 284 601
rect 285 600 286 601
rect 280 601 286 605
rect 280 605 281 606
rect 282 605 283 606
rect 283 605 284 606
rect 285 605 286 606
rect 680 940 681 941
rect 682 940 683 941
rect 683 940 684 941
rect 685 940 686 941
rect 680 941 686 945
rect 680 945 681 946
rect 682 945 683 946
rect 683 945 684 946
rect 685 945 686 946
rect 260 620 261 621
rect 262 620 263 621
rect 263 620 264 621
rect 265 620 266 621
rect 260 621 266 625
rect 260 625 261 626
rect 262 625 263 626
rect 263 625 264 626
rect 265 625 266 626
rect 700 540 701 541
rect 702 540 703 541
rect 703 540 704 541
rect 705 540 706 541
rect 700 541 706 545
rect 700 545 701 546
rect 702 545 703 546
rect 703 545 704 546
rect 705 545 706 546
rect 640 500 641 501
rect 642 500 643 501
rect 643 500 644 501
rect 645 500 646 501
rect 640 501 646 505
rect 640 505 641 506
rect 642 505 643 506
rect 643 505 644 506
rect 645 505 646 506
rect 900 700 901 701
rect 902 700 903 701
rect 903 700 904 701
rect 905 700 906 701
rect 900 701 906 705
rect 900 705 901 706
rect 902 705 903 706
rect 903 705 904 706
rect 905 705 906 706
rect 500 680 501 681
rect 502 680 503 681
rect 503 680 504 681
rect 505 680 506 681
rect 500 681 506 685
rect 500 685 501 686
rect 502 685 503 686
rect 503 685 504 686
rect 505 685 506 686
rect 480 940 481 941
rect 482 940 483 941
rect 483 940 484 941
rect 485 940 486 941
rect 480 941 486 945
rect 480 945 481 946
rect 482 945 483 946
rect 483 945 484 946
rect 485 945 486 946
rect 660 340 661 341
rect 662 340 663 341
rect 663 340 664 341
rect 665 340 666 341
rect 660 341 666 345
rect 660 345 661 346
rect 662 345 663 346
rect 663 345 664 346
rect 665 345 666 346
rect 440 740 441 741
rect 442 740 443 741
rect 443 740 444 741
rect 445 740 446 741
rect 440 741 446 745
rect 440 745 441 746
rect 442 745 443 746
rect 443 745 444 746
rect 445 745 446 746
rect 720 840 721 841
rect 722 840 723 841
rect 723 840 724 841
rect 725 840 726 841
rect 720 841 726 845
rect 720 845 721 846
rect 722 845 723 846
rect 723 845 724 846
rect 725 845 726 846
rect 700 860 701 861
rect 702 860 703 861
rect 703 860 704 861
rect 705 860 706 861
rect 700 861 706 865
rect 700 865 701 866
rect 702 865 703 866
rect 703 865 704 866
rect 705 865 706 866
rect 460 440 461 441
rect 462 440 463 441
rect 463 440 464 441
rect 465 440 466 441
rect 460 441 466 445
rect 460 445 461 446
rect 462 445 463 446
rect 463 445 464 446
rect 465 445 466 446
rect 740 340 741 341
rect 742 340 743 341
rect 743 340 744 341
rect 745 340 746 341
rect 740 341 746 345
rect 740 345 741 346
rect 742 345 743 346
rect 743 345 744 346
rect 745 345 746 346
rect 460 1040 461 1041
rect 462 1040 463 1041
rect 463 1040 464 1041
rect 465 1040 466 1041
rect 460 1041 466 1045
rect 460 1045 461 1046
rect 462 1045 463 1046
rect 463 1045 464 1046
rect 465 1045 466 1046
rect 640 300 641 301
rect 642 300 643 301
rect 643 300 644 301
rect 645 300 646 301
rect 640 301 646 305
rect 640 305 641 306
rect 642 305 643 306
rect 643 305 644 306
rect 645 305 646 306
rect 1040 660 1041 661
rect 1042 660 1043 661
rect 1043 660 1044 661
rect 1045 660 1046 661
rect 1040 661 1046 665
rect 1040 665 1041 666
rect 1042 665 1043 666
rect 1043 665 1044 666
rect 1045 665 1046 666
rect 500 420 501 421
rect 502 420 503 421
rect 503 420 504 421
rect 505 420 506 421
rect 500 421 506 425
rect 500 425 501 426
rect 502 425 503 426
rect 503 425 504 426
rect 505 425 506 426
rect 680 800 681 801
rect 682 800 683 801
rect 683 800 684 801
rect 685 800 686 801
rect 680 801 686 805
rect 680 805 681 806
rect 682 805 683 806
rect 683 805 684 806
rect 685 805 686 806
rect 720 620 721 621
rect 722 620 723 621
rect 723 620 724 621
rect 725 620 726 621
rect 720 621 726 625
rect 720 625 721 626
rect 722 625 723 626
rect 723 625 724 626
rect 725 625 726 626
rect 340 620 341 621
rect 342 620 343 621
rect 343 620 344 621
rect 345 620 346 621
rect 340 621 346 625
rect 340 625 341 626
rect 342 625 343 626
rect 343 625 344 626
rect 345 625 346 626
rect 420 640 421 641
rect 422 640 423 641
rect 423 640 424 641
rect 425 640 426 641
rect 420 641 426 645
rect 420 645 421 646
rect 422 645 423 646
rect 423 645 424 646
rect 425 645 426 646
rect 820 380 821 381
rect 822 380 823 381
rect 823 380 824 381
rect 825 380 826 381
rect 820 381 826 385
rect 820 385 821 386
rect 822 385 823 386
rect 823 385 824 386
rect 825 385 826 386
rect 360 520 361 521
rect 362 520 363 521
rect 363 520 364 521
rect 365 520 366 521
rect 360 521 366 525
rect 360 525 361 526
rect 362 525 363 526
rect 363 525 364 526
rect 365 525 366 526
rect 440 820 441 821
rect 442 820 443 821
rect 443 820 444 821
rect 445 820 446 821
rect 440 821 446 825
rect 440 825 441 826
rect 442 825 443 826
rect 443 825 444 826
rect 445 825 446 826
rect 560 920 561 921
rect 562 920 563 921
rect 563 920 564 921
rect 565 920 566 921
rect 560 921 566 925
rect 560 925 561 926
rect 562 925 563 926
rect 563 925 564 926
rect 565 925 566 926
rect 820 740 821 741
rect 822 740 823 741
rect 823 740 824 741
rect 825 740 826 741
rect 820 741 826 745
rect 820 745 821 746
rect 822 745 823 746
rect 823 745 824 746
rect 825 745 826 746
rect 920 760 921 761
rect 922 760 923 761
rect 923 760 924 761
rect 925 760 926 761
rect 920 761 926 765
rect 920 765 921 766
rect 922 765 923 766
rect 923 765 924 766
rect 925 765 926 766
rect 620 860 621 861
rect 622 860 623 861
rect 623 860 624 861
rect 625 860 626 861
rect 620 861 626 865
rect 620 865 621 866
rect 622 865 623 866
rect 623 865 624 866
rect 625 865 626 866
rect 680 380 681 381
rect 682 380 683 381
rect 683 380 684 381
rect 685 380 686 381
rect 680 381 686 385
rect 680 385 681 386
rect 682 385 683 386
rect 683 385 684 386
rect 685 385 686 386
rect 700 560 701 561
rect 702 560 703 561
rect 703 560 704 561
rect 705 560 706 561
rect 700 561 706 565
rect 700 565 701 566
rect 702 565 703 566
rect 703 565 704 566
rect 705 565 706 566
rect 920 500 921 501
rect 922 500 923 501
rect 923 500 924 501
rect 925 500 926 501
rect 920 501 926 505
rect 920 505 921 506
rect 922 505 923 506
rect 923 505 924 506
rect 925 505 926 506
rect 540 440 541 441
rect 542 440 543 441
rect 543 440 544 441
rect 545 440 546 441
rect 540 441 546 445
rect 540 445 541 446
rect 542 445 543 446
rect 543 445 544 446
rect 545 445 546 446
rect 500 540 501 541
rect 502 540 503 541
rect 503 540 504 541
rect 505 540 506 541
rect 500 541 506 545
rect 500 545 501 546
rect 502 545 503 546
rect 503 545 504 546
rect 505 545 506 546
rect 940 740 941 741
rect 942 740 943 741
rect 943 740 944 741
rect 945 740 946 741
rect 940 741 946 745
rect 940 745 941 746
rect 942 745 943 746
rect 943 745 944 746
rect 945 745 946 746
rect 840 860 841 861
rect 842 860 843 861
rect 843 860 844 861
rect 845 860 846 861
rect 840 861 846 865
rect 840 865 841 866
rect 842 865 843 866
rect 843 865 844 866
rect 845 865 846 866
rect 820 440 821 441
rect 822 440 823 441
rect 823 440 824 441
rect 825 440 826 441
rect 820 441 826 445
rect 820 445 821 446
rect 822 445 823 446
rect 823 445 824 446
rect 825 445 826 446
rect 940 640 941 641
rect 942 640 943 641
rect 943 640 944 641
rect 945 640 946 641
rect 940 641 946 645
rect 940 645 941 646
rect 942 645 943 646
rect 943 645 944 646
rect 945 645 946 646
rect 520 460 521 461
rect 522 460 523 461
rect 523 460 524 461
rect 525 460 526 461
rect 520 461 526 465
rect 520 465 521 466
rect 522 465 523 466
rect 523 465 524 466
rect 525 465 526 466
rect 1000 740 1001 741
rect 1002 740 1003 741
rect 1003 740 1004 741
rect 1005 740 1006 741
rect 1000 741 1006 745
rect 1000 745 1001 746
rect 1002 745 1003 746
rect 1003 745 1004 746
rect 1005 745 1006 746
rect 680 1000 681 1001
rect 682 1000 683 1001
rect 683 1000 684 1001
rect 685 1000 686 1001
rect 680 1001 686 1005
rect 680 1005 681 1006
rect 682 1005 683 1006
rect 683 1005 684 1006
rect 685 1005 686 1006
rect 500 640 501 641
rect 502 640 503 641
rect 503 640 504 641
rect 505 640 506 641
rect 500 641 506 645
rect 500 645 501 646
rect 502 645 503 646
rect 503 645 504 646
rect 505 645 506 646
rect 960 720 961 721
rect 962 720 963 721
rect 963 720 964 721
rect 965 720 966 721
rect 960 721 966 725
rect 960 725 961 726
rect 962 725 963 726
rect 963 725 964 726
rect 965 725 966 726
rect 700 600 701 601
rect 702 600 703 601
rect 703 600 704 601
rect 705 600 706 601
rect 700 601 706 605
rect 700 605 701 606
rect 702 605 703 606
rect 703 605 704 606
rect 705 605 706 606
rect 580 560 581 561
rect 582 560 583 561
rect 583 560 584 561
rect 585 560 586 561
rect 580 561 586 565
rect 580 565 581 566
rect 582 565 583 566
rect 583 565 584 566
rect 585 565 586 566
rect 760 900 761 901
rect 762 900 763 901
rect 763 900 764 901
rect 765 900 766 901
rect 760 901 766 905
rect 760 905 761 906
rect 762 905 763 906
rect 763 905 764 906
rect 765 905 766 906
rect 760 860 761 861
rect 762 860 763 861
rect 763 860 764 861
rect 765 860 766 861
rect 760 861 766 865
rect 760 865 761 866
rect 762 865 763 866
rect 763 865 764 866
rect 765 865 766 866
rect 600 660 601 661
rect 602 660 603 661
rect 603 660 604 661
rect 605 660 606 661
rect 600 661 606 665
rect 600 665 601 666
rect 602 665 603 666
rect 603 665 604 666
rect 605 665 606 666
rect 860 620 861 621
rect 862 620 863 621
rect 863 620 864 621
rect 865 620 866 621
rect 860 621 866 625
rect 860 625 861 626
rect 862 625 863 626
rect 863 625 864 626
rect 865 625 866 626
rect 900 500 901 501
rect 902 500 903 501
rect 903 500 904 501
rect 905 500 906 501
rect 900 501 906 505
rect 900 505 901 506
rect 902 505 903 506
rect 903 505 904 506
rect 905 505 906 506
rect 540 600 541 601
rect 542 600 543 601
rect 543 600 544 601
rect 545 600 546 601
rect 540 601 546 605
rect 540 605 541 606
rect 542 605 543 606
rect 543 605 544 606
rect 545 605 546 606
rect 680 420 681 421
rect 682 420 683 421
rect 683 420 684 421
rect 685 420 686 421
rect 680 421 686 425
rect 680 425 681 426
rect 682 425 683 426
rect 683 425 684 426
rect 685 425 686 426
rect 320 560 321 561
rect 322 560 323 561
rect 323 560 324 561
rect 325 560 326 561
rect 320 561 326 565
rect 320 565 321 566
rect 322 565 323 566
rect 323 565 324 566
rect 325 565 326 566
rect 560 900 561 901
rect 562 900 563 901
rect 563 900 564 901
rect 565 900 566 901
rect 560 901 566 905
rect 560 905 561 906
rect 562 905 563 906
rect 563 905 564 906
rect 565 905 566 906
rect 1020 680 1021 681
rect 1022 680 1023 681
rect 1023 680 1024 681
rect 1025 680 1026 681
rect 1020 681 1026 685
rect 1020 685 1021 686
rect 1022 685 1023 686
rect 1023 685 1024 686
rect 1025 685 1026 686
rect 480 600 481 601
rect 482 600 483 601
rect 483 600 484 601
rect 485 600 486 601
rect 480 601 486 605
rect 480 605 481 606
rect 482 605 483 606
rect 483 605 484 606
rect 485 605 486 606
rect 860 520 861 521
rect 862 520 863 521
rect 863 520 864 521
rect 865 520 866 521
rect 860 521 866 525
rect 860 525 861 526
rect 862 525 863 526
rect 863 525 864 526
rect 865 525 866 526
rect 740 780 741 781
rect 742 780 743 781
rect 743 780 744 781
rect 745 780 746 781
rect 740 781 746 785
rect 740 785 741 786
rect 742 785 743 786
rect 743 785 744 786
rect 745 785 746 786
rect 1040 700 1041 701
rect 1042 700 1043 701
rect 1043 700 1044 701
rect 1045 700 1046 701
rect 1040 701 1046 705
rect 1040 705 1041 706
rect 1042 705 1043 706
rect 1043 705 1044 706
rect 1045 705 1046 706
rect 880 720 881 721
rect 882 720 883 721
rect 883 720 884 721
rect 885 720 886 721
rect 880 721 886 725
rect 880 725 881 726
rect 882 725 883 726
rect 883 725 884 726
rect 885 725 886 726
rect 560 760 561 761
rect 562 760 563 761
rect 563 760 564 761
rect 565 760 566 761
rect 560 761 566 765
rect 560 765 561 766
rect 562 765 563 766
rect 563 765 564 766
rect 565 765 566 766
rect 820 500 821 501
rect 822 500 823 501
rect 823 500 824 501
rect 825 500 826 501
rect 820 501 826 505
rect 820 505 821 506
rect 822 505 823 506
rect 823 505 824 506
rect 825 505 826 506
rect 640 320 641 321
rect 642 320 643 321
rect 643 320 644 321
rect 645 320 646 321
rect 640 321 646 325
rect 640 325 641 326
rect 642 325 643 326
rect 643 325 644 326
rect 645 325 646 326
rect 760 800 761 801
rect 762 800 763 801
rect 763 800 764 801
rect 765 800 766 801
rect 760 801 766 805
rect 760 805 761 806
rect 762 805 763 806
rect 763 805 764 806
rect 765 805 766 806
rect 680 1040 681 1041
rect 682 1040 683 1041
rect 683 1040 684 1041
rect 685 1040 686 1041
rect 680 1041 686 1045
rect 680 1045 681 1046
rect 682 1045 683 1046
rect 683 1045 684 1046
rect 685 1045 686 1046
rect 640 920 641 921
rect 642 920 643 921
rect 643 920 644 921
rect 645 920 646 921
rect 640 921 646 925
rect 640 925 641 926
rect 642 925 643 926
rect 643 925 644 926
rect 645 925 646 926
rect 880 540 881 541
rect 882 540 883 541
rect 883 540 884 541
rect 885 540 886 541
rect 880 541 886 545
rect 880 545 881 546
rect 882 545 883 546
rect 883 545 884 546
rect 885 545 886 546
rect 620 800 621 801
rect 622 800 623 801
rect 623 800 624 801
rect 625 800 626 801
rect 620 801 626 805
rect 620 805 621 806
rect 622 805 623 806
rect 623 805 624 806
rect 625 805 626 806
rect 380 520 381 521
rect 382 520 383 521
rect 383 520 384 521
rect 385 520 386 521
rect 380 521 386 525
rect 380 525 381 526
rect 382 525 383 526
rect 383 525 384 526
rect 385 525 386 526
rect 580 620 581 621
rect 582 620 583 621
rect 583 620 584 621
rect 585 620 586 621
rect 580 621 586 625
rect 580 625 581 626
rect 582 625 583 626
rect 583 625 584 626
rect 585 625 586 626
rect 960 600 961 601
rect 962 600 963 601
rect 963 600 964 601
rect 965 600 966 601
rect 960 601 966 605
rect 960 605 961 606
rect 962 605 963 606
rect 963 605 964 606
rect 965 605 966 606
rect 740 480 741 481
rect 742 480 743 481
rect 743 480 744 481
rect 745 480 746 481
rect 740 481 746 485
rect 740 485 741 486
rect 742 485 743 486
rect 743 485 744 486
rect 745 485 746 486
rect 800 580 801 581
rect 802 580 803 581
rect 803 580 804 581
rect 805 580 806 581
rect 800 581 806 585
rect 800 585 801 586
rect 802 585 803 586
rect 803 585 804 586
rect 805 585 806 586
rect 420 460 421 461
rect 422 460 423 461
rect 423 460 424 461
rect 425 460 426 461
rect 420 461 426 465
rect 420 465 421 466
rect 422 465 423 466
rect 423 465 424 466
rect 425 465 426 466
rect 500 460 501 461
rect 502 460 503 461
rect 503 460 504 461
rect 505 460 506 461
rect 500 461 506 465
rect 500 465 501 466
rect 502 465 503 466
rect 503 465 504 466
rect 505 465 506 466
rect 720 780 721 781
rect 722 780 723 781
rect 723 780 724 781
rect 725 780 726 781
rect 720 781 726 785
rect 720 785 721 786
rect 722 785 723 786
rect 723 785 724 786
rect 725 785 726 786
rect 580 940 581 941
rect 582 940 583 941
rect 583 940 584 941
rect 585 940 586 941
rect 580 941 586 945
rect 580 945 581 946
rect 582 945 583 946
rect 583 945 584 946
rect 585 945 586 946
rect 640 380 641 381
rect 642 380 643 381
rect 643 380 644 381
rect 645 380 646 381
rect 640 381 646 385
rect 640 385 641 386
rect 642 385 643 386
rect 643 385 644 386
rect 645 385 646 386
rect 900 640 901 641
rect 902 640 903 641
rect 903 640 904 641
rect 905 640 906 641
rect 900 641 906 645
rect 900 645 901 646
rect 902 645 903 646
rect 903 645 904 646
rect 905 645 906 646
rect 780 820 781 821
rect 782 820 783 821
rect 783 820 784 821
rect 785 820 786 821
rect 780 821 786 825
rect 780 825 781 826
rect 782 825 783 826
rect 783 825 784 826
rect 785 825 786 826
rect 340 820 341 821
rect 342 820 343 821
rect 343 820 344 821
rect 345 820 346 821
rect 340 821 346 825
rect 340 825 341 826
rect 342 825 343 826
rect 343 825 344 826
rect 345 825 346 826
rect 620 280 621 281
rect 622 280 623 281
rect 623 280 624 281
rect 625 280 626 281
rect 620 281 626 285
rect 620 285 621 286
rect 622 285 623 286
rect 623 285 624 286
rect 625 285 626 286
rect 580 360 581 361
rect 582 360 583 361
rect 583 360 584 361
rect 585 360 586 361
rect 580 361 586 365
rect 580 365 581 366
rect 582 365 583 366
rect 583 365 584 366
rect 585 365 586 366
rect 800 740 801 741
rect 802 740 803 741
rect 803 740 804 741
rect 805 740 806 741
rect 800 741 806 745
rect 800 745 801 746
rect 802 745 803 746
rect 803 745 804 746
rect 805 745 806 746
rect 740 820 741 821
rect 742 820 743 821
rect 743 820 744 821
rect 745 820 746 821
rect 740 821 746 825
rect 740 825 741 826
rect 742 825 743 826
rect 743 825 744 826
rect 745 825 746 826
rect 240 700 241 701
rect 242 700 243 701
rect 243 700 244 701
rect 245 700 246 701
rect 240 701 246 705
rect 240 705 241 706
rect 242 705 243 706
rect 243 705 244 706
rect 245 705 246 706
rect 460 680 461 681
rect 462 680 463 681
rect 463 680 464 681
rect 465 680 466 681
rect 460 681 466 685
rect 460 685 461 686
rect 462 685 463 686
rect 463 685 464 686
rect 465 685 466 686
rect 940 700 941 701
rect 942 700 943 701
rect 943 700 944 701
rect 945 700 946 701
rect 940 701 946 705
rect 940 705 941 706
rect 942 705 943 706
rect 943 705 944 706
rect 945 705 946 706
rect 760 920 761 921
rect 762 920 763 921
rect 763 920 764 921
rect 765 920 766 921
rect 760 921 766 925
rect 760 925 761 926
rect 762 925 763 926
rect 763 925 764 926
rect 765 925 766 926
rect 800 840 801 841
rect 802 840 803 841
rect 803 840 804 841
rect 805 840 806 841
rect 800 841 806 845
rect 800 845 801 846
rect 802 845 803 846
rect 803 845 804 846
rect 805 845 806 846
rect 600 360 601 361
rect 602 360 603 361
rect 603 360 604 361
rect 605 360 606 361
rect 600 361 606 365
rect 600 365 601 366
rect 602 365 603 366
rect 603 365 604 366
rect 605 365 606 366
rect 820 520 821 521
rect 822 520 823 521
rect 823 520 824 521
rect 825 520 826 521
rect 820 521 826 525
rect 820 525 821 526
rect 822 525 823 526
rect 823 525 824 526
rect 825 525 826 526
rect 840 800 841 801
rect 842 800 843 801
rect 843 800 844 801
rect 845 800 846 801
rect 840 801 846 805
rect 840 805 841 806
rect 842 805 843 806
rect 843 805 844 806
rect 845 805 846 806
rect 520 720 521 721
rect 522 720 523 721
rect 523 720 524 721
rect 525 720 526 721
rect 520 721 526 725
rect 520 725 521 726
rect 522 725 523 726
rect 523 725 524 726
rect 525 725 526 726
rect 360 620 361 621
rect 362 620 363 621
rect 363 620 364 621
rect 365 620 366 621
rect 360 621 366 625
rect 360 625 361 626
rect 362 625 363 626
rect 363 625 364 626
rect 365 625 366 626
rect 700 640 701 641
rect 702 640 703 641
rect 703 640 704 641
rect 705 640 706 641
rect 700 641 706 645
rect 700 645 701 646
rect 702 645 703 646
rect 703 645 704 646
rect 705 645 706 646
rect 460 840 461 841
rect 462 840 463 841
rect 463 840 464 841
rect 465 840 466 841
rect 460 841 466 845
rect 460 845 461 846
rect 462 845 463 846
rect 463 845 464 846
rect 465 845 466 846
rect 360 660 361 661
rect 362 660 363 661
rect 363 660 364 661
rect 365 660 366 661
rect 360 661 366 665
rect 360 665 361 666
rect 362 665 363 666
rect 363 665 364 666
rect 365 665 366 666
rect 720 320 721 321
rect 722 320 723 321
rect 723 320 724 321
rect 725 320 726 321
rect 720 321 726 325
rect 720 325 721 326
rect 722 325 723 326
rect 723 325 724 326
rect 725 325 726 326
rect 340 640 341 641
rect 342 640 343 641
rect 343 640 344 641
rect 345 640 346 641
rect 340 641 346 645
rect 340 645 341 646
rect 342 645 343 646
rect 343 645 344 646
rect 345 645 346 646
rect 400 680 401 681
rect 402 680 403 681
rect 403 680 404 681
rect 405 680 406 681
rect 400 681 406 685
rect 400 685 401 686
rect 402 685 403 686
rect 403 685 404 686
rect 405 685 406 686
rect 980 580 981 581
rect 982 580 983 581
rect 983 580 984 581
rect 985 580 986 581
rect 980 581 986 585
rect 980 585 981 586
rect 982 585 983 586
rect 983 585 984 586
rect 985 585 986 586
rect 560 1020 561 1021
rect 562 1020 563 1021
rect 563 1020 564 1021
rect 565 1020 566 1021
rect 560 1021 566 1025
rect 560 1025 561 1026
rect 562 1025 563 1026
rect 563 1025 564 1026
rect 565 1025 566 1026
rect 780 420 781 421
rect 782 420 783 421
rect 783 420 784 421
rect 785 420 786 421
rect 780 421 786 425
rect 780 425 781 426
rect 782 425 783 426
rect 783 425 784 426
rect 785 425 786 426
rect 800 400 801 401
rect 802 400 803 401
rect 803 400 804 401
rect 805 400 806 401
rect 800 401 806 405
rect 800 405 801 406
rect 802 405 803 406
rect 803 405 804 406
rect 805 405 806 406
rect 660 380 661 381
rect 662 380 663 381
rect 663 380 664 381
rect 665 380 666 381
rect 660 381 666 385
rect 660 385 661 386
rect 662 385 663 386
rect 663 385 664 386
rect 665 385 666 386
rect 400 540 401 541
rect 402 540 403 541
rect 403 540 404 541
rect 405 540 406 541
rect 400 541 406 545
rect 400 545 401 546
rect 402 545 403 546
rect 403 545 404 546
rect 405 545 406 546
rect 400 520 401 521
rect 402 520 403 521
rect 403 520 404 521
rect 405 520 406 521
rect 400 521 406 525
rect 400 525 401 526
rect 402 525 403 526
rect 403 525 404 526
rect 405 525 406 526
rect 420 700 421 701
rect 422 700 423 701
rect 423 700 424 701
rect 425 700 426 701
rect 420 701 426 705
rect 420 705 421 706
rect 422 705 423 706
rect 423 705 424 706
rect 425 705 426 706
rect 860 900 861 901
rect 862 900 863 901
rect 863 900 864 901
rect 865 900 866 901
rect 860 901 866 905
rect 860 905 861 906
rect 862 905 863 906
rect 863 905 864 906
rect 865 905 866 906
rect 520 880 521 881
rect 522 880 523 881
rect 523 880 524 881
rect 525 880 526 881
rect 520 881 526 885
rect 520 885 521 886
rect 522 885 523 886
rect 523 885 524 886
rect 525 885 526 886
rect 820 680 821 681
rect 822 680 823 681
rect 823 680 824 681
rect 825 680 826 681
rect 820 681 826 685
rect 820 685 821 686
rect 822 685 823 686
rect 823 685 824 686
rect 825 685 826 686
rect 860 880 861 881
rect 862 880 863 881
rect 863 880 864 881
rect 865 880 866 881
rect 860 881 866 885
rect 860 885 861 886
rect 862 885 863 886
rect 863 885 864 886
rect 865 885 866 886
rect 940 800 941 801
rect 942 800 943 801
rect 943 800 944 801
rect 945 800 946 801
rect 940 801 946 805
rect 940 805 941 806
rect 942 805 943 806
rect 943 805 944 806
rect 945 805 946 806
rect 580 980 581 981
rect 582 980 583 981
rect 583 980 584 981
rect 585 980 586 981
rect 580 981 586 985
rect 580 985 581 986
rect 582 985 583 986
rect 583 985 584 986
rect 585 985 586 986
rect 620 360 621 361
rect 622 360 623 361
rect 623 360 624 361
rect 625 360 626 361
rect 620 361 626 365
rect 620 365 621 366
rect 622 365 623 366
rect 623 365 624 366
rect 625 365 626 366
rect 980 660 981 661
rect 982 660 983 661
rect 983 660 984 661
rect 985 660 986 661
rect 980 661 986 665
rect 980 665 981 666
rect 982 665 983 666
rect 983 665 984 666
rect 985 665 986 666
rect 860 860 861 861
rect 862 860 863 861
rect 863 860 864 861
rect 865 860 866 861
rect 860 861 866 865
rect 860 865 861 866
rect 862 865 863 866
rect 863 865 864 866
rect 865 865 866 866
rect 660 940 661 941
rect 662 940 663 941
rect 663 940 664 941
rect 665 940 666 941
rect 660 941 666 945
rect 660 945 661 946
rect 662 945 663 946
rect 663 945 664 946
rect 665 945 666 946
rect 720 880 721 881
rect 722 880 723 881
rect 723 880 724 881
rect 725 880 726 881
rect 720 881 726 885
rect 720 885 721 886
rect 722 885 723 886
rect 723 885 724 886
rect 725 885 726 886
rect 820 800 821 801
rect 822 800 823 801
rect 823 800 824 801
rect 825 800 826 801
rect 820 801 826 805
rect 820 805 821 806
rect 822 805 823 806
rect 823 805 824 806
rect 825 805 826 806
rect 760 980 761 981
rect 762 980 763 981
rect 763 980 764 981
rect 765 980 766 981
rect 760 981 766 985
rect 760 985 761 986
rect 762 985 763 986
rect 763 985 764 986
rect 765 985 766 986
rect 800 360 801 361
rect 802 360 803 361
rect 803 360 804 361
rect 805 360 806 361
rect 800 361 806 365
rect 800 365 801 366
rect 802 365 803 366
rect 803 365 804 366
rect 805 365 806 366
rect 380 680 381 681
rect 382 680 383 681
rect 383 680 384 681
rect 385 680 386 681
rect 380 681 386 685
rect 380 685 381 686
rect 382 685 383 686
rect 383 685 384 686
rect 385 685 386 686
rect 340 720 341 721
rect 342 720 343 721
rect 343 720 344 721
rect 345 720 346 721
rect 340 721 346 725
rect 340 725 341 726
rect 342 725 343 726
rect 343 725 344 726
rect 345 725 346 726
rect 700 920 701 921
rect 702 920 703 921
rect 703 920 704 921
rect 705 920 706 921
rect 700 921 706 925
rect 700 925 701 926
rect 702 925 703 926
rect 703 925 704 926
rect 705 925 706 926
rect 740 420 741 421
rect 742 420 743 421
rect 743 420 744 421
rect 745 420 746 421
rect 740 421 746 425
rect 740 425 741 426
rect 742 425 743 426
rect 743 425 744 426
rect 745 425 746 426
rect 760 960 761 961
rect 762 960 763 961
rect 763 960 764 961
rect 765 960 766 961
rect 760 961 766 965
rect 760 965 761 966
rect 762 965 763 966
rect 763 965 764 966
rect 765 965 766 966
rect 780 780 781 781
rect 782 780 783 781
rect 783 780 784 781
rect 785 780 786 781
rect 780 781 786 785
rect 780 785 781 786
rect 782 785 783 786
rect 783 785 784 786
rect 785 785 786 786
rect 900 760 901 761
rect 902 760 903 761
rect 903 760 904 761
rect 905 760 906 761
rect 900 761 906 765
rect 900 765 901 766
rect 902 765 903 766
rect 903 765 904 766
rect 905 765 906 766
rect 660 1080 661 1081
rect 662 1080 663 1081
rect 663 1080 664 1081
rect 665 1080 666 1081
rect 660 1081 666 1085
rect 660 1085 661 1086
rect 662 1085 663 1086
rect 663 1085 664 1086
rect 665 1085 666 1086
rect 600 1020 601 1021
rect 602 1020 603 1021
rect 603 1020 604 1021
rect 605 1020 606 1021
rect 600 1021 606 1025
rect 600 1025 601 1026
rect 602 1025 603 1026
rect 603 1025 604 1026
rect 605 1025 606 1026
rect 480 560 481 561
rect 482 560 483 561
rect 483 560 484 561
rect 485 560 486 561
rect 480 561 486 565
rect 480 565 481 566
rect 482 565 483 566
rect 483 565 484 566
rect 485 565 486 566
rect 540 920 541 921
rect 542 920 543 921
rect 543 920 544 921
rect 545 920 546 921
rect 540 921 546 925
rect 540 925 541 926
rect 542 925 543 926
rect 543 925 544 926
rect 545 925 546 926
rect 720 560 721 561
rect 722 560 723 561
rect 723 560 724 561
rect 725 560 726 561
rect 720 561 726 565
rect 720 565 721 566
rect 722 565 723 566
rect 723 565 724 566
rect 725 565 726 566
rect 780 480 781 481
rect 782 480 783 481
rect 783 480 784 481
rect 785 480 786 481
rect 780 481 786 485
rect 780 485 781 486
rect 782 485 783 486
rect 783 485 784 486
rect 785 485 786 486
rect 940 780 941 781
rect 942 780 943 781
rect 943 780 944 781
rect 945 780 946 781
rect 940 781 946 785
rect 940 785 941 786
rect 942 785 943 786
rect 943 785 944 786
rect 945 785 946 786
rect 1000 620 1001 621
rect 1002 620 1003 621
rect 1003 620 1004 621
rect 1005 620 1006 621
rect 1000 621 1006 625
rect 1000 625 1001 626
rect 1002 625 1003 626
rect 1003 625 1004 626
rect 1005 625 1006 626
rect 620 440 621 441
rect 622 440 623 441
rect 623 440 624 441
rect 625 440 626 441
rect 620 441 626 445
rect 620 445 621 446
rect 622 445 623 446
rect 623 445 624 446
rect 625 445 626 446
rect 620 900 621 901
rect 622 900 623 901
rect 623 900 624 901
rect 625 900 626 901
rect 620 901 626 905
rect 620 905 621 906
rect 622 905 623 906
rect 623 905 624 906
rect 625 905 626 906
rect 280 720 281 721
rect 282 720 283 721
rect 283 720 284 721
rect 285 720 286 721
rect 280 721 286 725
rect 280 725 281 726
rect 282 725 283 726
rect 283 725 284 726
rect 285 725 286 726
rect 920 640 921 641
rect 922 640 923 641
rect 923 640 924 641
rect 925 640 926 641
rect 920 641 926 645
rect 920 645 921 646
rect 922 645 923 646
rect 923 645 924 646
rect 925 645 926 646
rect 720 400 721 401
rect 722 400 723 401
rect 723 400 724 401
rect 725 400 726 401
rect 720 401 726 405
rect 720 405 721 406
rect 722 405 723 406
rect 723 405 724 406
rect 725 405 726 406
rect 380 800 381 801
rect 382 800 383 801
rect 383 800 384 801
rect 385 800 386 801
rect 380 801 386 805
rect 380 805 381 806
rect 382 805 383 806
rect 383 805 384 806
rect 385 805 386 806
rect 860 480 861 481
rect 862 480 863 481
rect 863 480 864 481
rect 865 480 866 481
rect 860 481 866 485
rect 860 485 861 486
rect 862 485 863 486
rect 863 485 864 486
rect 865 485 866 486
rect 780 600 781 601
rect 782 600 783 601
rect 783 600 784 601
rect 785 600 786 601
rect 780 601 786 605
rect 780 605 781 606
rect 782 605 783 606
rect 783 605 784 606
rect 785 605 786 606
rect 640 580 641 581
rect 642 580 643 581
rect 643 580 644 581
rect 645 580 646 581
rect 640 581 646 585
rect 640 585 641 586
rect 642 585 643 586
rect 643 585 644 586
rect 645 585 646 586
rect 340 600 341 601
rect 342 600 343 601
rect 343 600 344 601
rect 345 600 346 601
rect 340 601 346 605
rect 340 605 341 606
rect 342 605 343 606
rect 343 605 344 606
rect 345 605 346 606
rect 920 540 921 541
rect 922 540 923 541
rect 923 540 924 541
rect 925 540 926 541
rect 920 541 926 545
rect 920 545 921 546
rect 922 545 923 546
rect 923 545 924 546
rect 925 545 926 546
rect 780 380 781 381
rect 782 380 783 381
rect 783 380 784 381
rect 785 380 786 381
rect 780 381 786 385
rect 780 385 781 386
rect 782 385 783 386
rect 783 385 784 386
rect 785 385 786 386
rect 520 960 521 961
rect 522 960 523 961
rect 523 960 524 961
rect 525 960 526 961
rect 520 961 526 965
rect 520 965 521 966
rect 522 965 523 966
rect 523 965 524 966
rect 525 965 526 966
rect 1020 600 1021 601
rect 1022 600 1023 601
rect 1023 600 1024 601
rect 1025 600 1026 601
rect 1020 601 1026 605
rect 1020 605 1021 606
rect 1022 605 1023 606
rect 1023 605 1024 606
rect 1025 605 1026 606
rect 720 340 721 341
rect 722 340 723 341
rect 723 340 724 341
rect 725 340 726 341
rect 720 341 726 345
rect 720 345 721 346
rect 722 345 723 346
rect 723 345 724 346
rect 725 345 726 346
rect 480 860 481 861
rect 482 860 483 861
rect 483 860 484 861
rect 485 860 486 861
rect 480 861 486 865
rect 480 865 481 866
rect 482 865 483 866
rect 483 865 484 866
rect 485 865 486 866
rect 360 680 361 681
rect 362 680 363 681
rect 363 680 364 681
rect 365 680 366 681
rect 360 681 366 685
rect 360 685 361 686
rect 362 685 363 686
rect 363 685 364 686
rect 365 685 366 686
rect 300 600 301 601
rect 302 600 303 601
rect 303 600 304 601
rect 305 600 306 601
rect 300 601 306 605
rect 300 605 301 606
rect 302 605 303 606
rect 303 605 304 606
rect 305 605 306 606
rect 700 340 701 341
rect 702 340 703 341
rect 703 340 704 341
rect 705 340 706 341
rect 700 341 706 345
rect 700 345 701 346
rect 702 345 703 346
rect 703 345 704 346
rect 705 345 706 346
rect 640 980 641 981
rect 642 980 643 981
rect 643 980 644 981
rect 645 980 646 981
rect 640 981 646 985
rect 640 985 641 986
rect 642 985 643 986
rect 643 985 644 986
rect 645 985 646 986
rect 360 760 361 761
rect 362 760 363 761
rect 363 760 364 761
rect 365 760 366 761
rect 360 761 366 765
rect 360 765 361 766
rect 362 765 363 766
rect 363 765 364 766
rect 365 765 366 766
rect 380 780 381 781
rect 382 780 383 781
rect 383 780 384 781
rect 385 780 386 781
rect 380 781 386 785
rect 380 785 381 786
rect 382 785 383 786
rect 383 785 384 786
rect 385 785 386 786
rect 900 680 901 681
rect 902 680 903 681
rect 903 680 904 681
rect 905 680 906 681
rect 900 681 906 685
rect 900 685 901 686
rect 902 685 903 686
rect 903 685 904 686
rect 905 685 906 686
rect 780 660 781 661
rect 782 660 783 661
rect 783 660 784 661
rect 785 660 786 661
rect 780 661 786 665
rect 780 665 781 666
rect 782 665 783 666
rect 783 665 784 666
rect 785 665 786 666
rect 800 680 801 681
rect 802 680 803 681
rect 803 680 804 681
rect 805 680 806 681
rect 800 681 806 685
rect 800 685 801 686
rect 802 685 803 686
rect 803 685 804 686
rect 805 685 806 686
rect 680 720 681 721
rect 682 720 683 721
rect 683 720 684 721
rect 685 720 686 721
rect 680 721 686 725
rect 680 725 681 726
rect 682 725 683 726
rect 683 725 684 726
rect 685 725 686 726
rect 500 740 501 741
rect 502 740 503 741
rect 503 740 504 741
rect 505 740 506 741
rect 500 741 506 745
rect 500 745 501 746
rect 502 745 503 746
rect 503 745 504 746
rect 505 745 506 746
rect 720 580 721 581
rect 722 580 723 581
rect 723 580 724 581
rect 725 580 726 581
rect 720 581 726 585
rect 720 585 721 586
rect 722 585 723 586
rect 723 585 724 586
rect 725 585 726 586
rect 280 700 281 701
rect 282 700 283 701
rect 283 700 284 701
rect 285 700 286 701
rect 280 701 286 705
rect 280 705 281 706
rect 282 705 283 706
rect 283 705 284 706
rect 285 705 286 706
rect 840 560 841 561
rect 842 560 843 561
rect 843 560 844 561
rect 845 560 846 561
rect 840 561 846 565
rect 840 565 841 566
rect 842 565 843 566
rect 843 565 844 566
rect 845 565 846 566
rect 380 760 381 761
rect 382 760 383 761
rect 383 760 384 761
rect 385 760 386 761
rect 380 761 386 765
rect 380 765 381 766
rect 382 765 383 766
rect 383 765 384 766
rect 385 765 386 766
rect 620 640 621 641
rect 622 640 623 641
rect 623 640 624 641
rect 625 640 626 641
rect 620 641 626 645
rect 620 645 621 646
rect 622 645 623 646
rect 623 645 624 646
rect 625 645 626 646
rect 540 880 541 881
rect 542 880 543 881
rect 543 880 544 881
rect 545 880 546 881
rect 540 881 546 885
rect 540 885 541 886
rect 542 885 543 886
rect 543 885 544 886
rect 545 885 546 886
rect 1020 620 1021 621
rect 1022 620 1023 621
rect 1023 620 1024 621
rect 1025 620 1026 621
rect 1020 621 1026 625
rect 1020 625 1021 626
rect 1022 625 1023 626
rect 1023 625 1024 626
rect 1025 625 1026 626
rect 780 560 781 561
rect 782 560 783 561
rect 783 560 784 561
rect 785 560 786 561
rect 780 561 786 565
rect 780 565 781 566
rect 782 565 783 566
rect 783 565 784 566
rect 785 565 786 566
rect 460 660 461 661
rect 462 660 463 661
rect 463 660 464 661
rect 465 660 466 661
rect 460 661 466 665
rect 460 665 461 666
rect 462 665 463 666
rect 463 665 464 666
rect 465 665 466 666
rect 760 540 761 541
rect 762 540 763 541
rect 763 540 764 541
rect 765 540 766 541
rect 760 541 766 545
rect 760 545 761 546
rect 762 545 763 546
rect 763 545 764 546
rect 765 545 766 546
rect 420 720 421 721
rect 422 720 423 721
rect 423 720 424 721
rect 425 720 426 721
rect 420 721 426 725
rect 420 725 421 726
rect 422 725 423 726
rect 423 725 424 726
rect 425 725 426 726
rect 540 520 541 521
rect 542 520 543 521
rect 543 520 544 521
rect 545 520 546 521
rect 540 521 546 525
rect 540 525 541 526
rect 542 525 543 526
rect 543 525 544 526
rect 545 525 546 526
rect 520 820 521 821
rect 522 820 523 821
rect 523 820 524 821
rect 525 820 526 821
rect 520 821 526 825
rect 520 825 521 826
rect 522 825 523 826
rect 523 825 524 826
rect 525 825 526 826
rect 960 560 961 561
rect 962 560 963 561
rect 963 560 964 561
rect 965 560 966 561
rect 960 561 966 565
rect 960 565 961 566
rect 962 565 963 566
rect 963 565 964 566
rect 965 565 966 566
rect 580 580 581 581
rect 582 580 583 581
rect 583 580 584 581
rect 585 580 586 581
rect 580 581 586 585
rect 580 585 581 586
rect 582 585 583 586
rect 583 585 584 586
rect 585 585 586 586
rect 800 760 801 761
rect 802 760 803 761
rect 803 760 804 761
rect 805 760 806 761
rect 800 761 806 765
rect 800 765 801 766
rect 802 765 803 766
rect 803 765 804 766
rect 805 765 806 766
rect 880 560 881 561
rect 882 560 883 561
rect 883 560 884 561
rect 885 560 886 561
rect 880 561 886 565
rect 880 565 881 566
rect 882 565 883 566
rect 883 565 884 566
rect 885 565 886 566
rect 760 580 761 581
rect 762 580 763 581
rect 763 580 764 581
rect 765 580 766 581
rect 760 581 766 585
rect 760 585 761 586
rect 762 585 763 586
rect 763 585 764 586
rect 765 585 766 586
rect 740 840 741 841
rect 742 840 743 841
rect 743 840 744 841
rect 745 840 746 841
rect 740 841 746 845
rect 740 845 741 846
rect 742 845 743 846
rect 743 845 744 846
rect 745 845 746 846
rect 640 600 641 601
rect 642 600 643 601
rect 643 600 644 601
rect 645 600 646 601
rect 640 601 646 605
rect 640 605 641 606
rect 642 605 643 606
rect 643 605 644 606
rect 645 605 646 606
rect 780 740 781 741
rect 782 740 783 741
rect 783 740 784 741
rect 785 740 786 741
rect 780 741 786 745
rect 780 745 781 746
rect 782 745 783 746
rect 783 745 784 746
rect 785 745 786 746
rect 780 720 781 721
rect 782 720 783 721
rect 783 720 784 721
rect 785 720 786 721
rect 780 721 786 725
rect 780 725 781 726
rect 782 725 783 726
rect 783 725 784 726
rect 785 725 786 726
rect 600 700 601 701
rect 602 700 603 701
rect 603 700 604 701
rect 605 700 606 701
rect 600 701 606 705
rect 600 705 601 706
rect 602 705 603 706
rect 603 705 604 706
rect 605 705 606 706
rect 980 740 981 741
rect 982 740 983 741
rect 983 740 984 741
rect 985 740 986 741
rect 980 741 986 745
rect 980 745 981 746
rect 982 745 983 746
rect 983 745 984 746
rect 985 745 986 746
rect 320 800 321 801
rect 322 800 323 801
rect 323 800 324 801
rect 325 800 326 801
rect 320 801 326 805
rect 320 805 321 806
rect 322 805 323 806
rect 323 805 324 806
rect 325 805 326 806
rect 900 600 901 601
rect 902 600 903 601
rect 903 600 904 601
rect 905 600 906 601
rect 900 601 906 605
rect 900 605 901 606
rect 902 605 903 606
rect 903 605 904 606
rect 905 605 906 606
rect 1000 720 1001 721
rect 1002 720 1003 721
rect 1003 720 1004 721
rect 1005 720 1006 721
rect 1000 721 1006 725
rect 1000 725 1001 726
rect 1002 725 1003 726
rect 1003 725 1004 726
rect 1005 725 1006 726
rect 580 880 581 881
rect 582 880 583 881
rect 583 880 584 881
rect 585 880 586 881
rect 580 881 586 885
rect 580 885 581 886
rect 582 885 583 886
rect 583 885 584 886
rect 585 885 586 886
rect 620 460 621 461
rect 622 460 623 461
rect 623 460 624 461
rect 625 460 626 461
rect 620 461 626 465
rect 620 465 621 466
rect 622 465 623 466
rect 623 465 624 466
rect 625 465 626 466
rect 840 440 841 441
rect 842 440 843 441
rect 843 440 844 441
rect 845 440 846 441
rect 840 441 846 445
rect 840 445 841 446
rect 842 445 843 446
rect 843 445 844 446
rect 845 445 846 446
rect 800 780 801 781
rect 802 780 803 781
rect 803 780 804 781
rect 805 780 806 781
rect 800 781 806 785
rect 800 785 801 786
rect 802 785 803 786
rect 803 785 804 786
rect 805 785 806 786
rect 640 880 641 881
rect 642 880 643 881
rect 643 880 644 881
rect 645 880 646 881
rect 640 881 646 885
rect 640 885 641 886
rect 642 885 643 886
rect 643 885 644 886
rect 645 885 646 886
rect 840 920 841 921
rect 842 920 843 921
rect 843 920 844 921
rect 845 920 846 921
rect 840 921 846 925
rect 840 925 841 926
rect 842 925 843 926
rect 843 925 844 926
rect 845 925 846 926
rect 700 380 701 381
rect 702 380 703 381
rect 703 380 704 381
rect 705 380 706 381
rect 700 381 706 385
rect 700 385 701 386
rect 702 385 703 386
rect 703 385 704 386
rect 705 385 706 386
rect 600 620 601 621
rect 602 620 603 621
rect 603 620 604 621
rect 605 620 606 621
rect 600 621 606 625
rect 600 625 601 626
rect 602 625 603 626
rect 603 625 604 626
rect 605 625 606 626
rect 540 660 541 661
rect 542 660 543 661
rect 543 660 544 661
rect 545 660 546 661
rect 540 661 546 665
rect 540 665 541 666
rect 542 665 543 666
rect 543 665 544 666
rect 545 665 546 666
rect 640 1060 641 1061
rect 642 1060 643 1061
rect 643 1060 644 1061
rect 645 1060 646 1061
rect 640 1061 646 1065
rect 640 1065 641 1066
rect 642 1065 643 1066
rect 643 1065 644 1066
rect 645 1065 646 1066
rect 380 820 381 821
rect 382 820 383 821
rect 383 820 384 821
rect 385 820 386 821
rect 380 821 386 825
rect 380 825 381 826
rect 382 825 383 826
rect 383 825 384 826
rect 385 825 386 826
rect 620 1080 621 1081
rect 622 1080 623 1081
rect 623 1080 624 1081
rect 625 1080 626 1081
rect 620 1081 626 1085
rect 620 1085 621 1086
rect 622 1085 623 1086
rect 623 1085 624 1086
rect 625 1085 626 1086
rect 780 960 781 961
rect 782 960 783 961
rect 783 960 784 961
rect 785 960 786 961
rect 780 961 786 965
rect 780 965 781 966
rect 782 965 783 966
rect 783 965 784 966
rect 785 965 786 966
rect 660 300 661 301
rect 662 300 663 301
rect 663 300 664 301
rect 665 300 666 301
rect 660 301 666 305
rect 660 305 661 306
rect 662 305 663 306
rect 663 305 664 306
rect 665 305 666 306
rect 520 440 521 441
rect 522 440 523 441
rect 523 440 524 441
rect 525 440 526 441
rect 520 441 526 445
rect 520 445 521 446
rect 522 445 523 446
rect 523 445 524 446
rect 525 445 526 446
rect 800 440 801 441
rect 802 440 803 441
rect 803 440 804 441
rect 805 440 806 441
rect 800 441 806 445
rect 800 445 801 446
rect 802 445 803 446
rect 803 445 804 446
rect 805 445 806 446
rect 340 780 341 781
rect 342 780 343 781
rect 343 780 344 781
rect 345 780 346 781
rect 340 781 346 785
rect 340 785 341 786
rect 342 785 343 786
rect 343 785 344 786
rect 345 785 346 786
rect 540 500 541 501
rect 542 500 543 501
rect 543 500 544 501
rect 545 500 546 501
rect 540 501 546 505
rect 540 505 541 506
rect 542 505 543 506
rect 543 505 544 506
rect 545 505 546 506
rect 560 700 561 701
rect 562 700 563 701
rect 563 700 564 701
rect 565 700 566 701
rect 560 701 566 705
rect 560 705 561 706
rect 562 705 563 706
rect 563 705 564 706
rect 565 705 566 706
rect 440 580 441 581
rect 442 580 443 581
rect 443 580 444 581
rect 445 580 446 581
rect 440 581 446 585
rect 440 585 441 586
rect 442 585 443 586
rect 443 585 444 586
rect 445 585 446 586
rect 540 980 541 981
rect 542 980 543 981
rect 543 980 544 981
rect 545 980 546 981
rect 540 981 546 985
rect 540 985 541 986
rect 542 985 543 986
rect 543 985 544 986
rect 545 985 546 986
rect 420 620 421 621
rect 422 620 423 621
rect 423 620 424 621
rect 425 620 426 621
rect 420 621 426 625
rect 420 625 421 626
rect 422 625 423 626
rect 423 625 424 626
rect 425 625 426 626
rect 300 700 301 701
rect 302 700 303 701
rect 303 700 304 701
rect 305 700 306 701
rect 300 701 306 705
rect 300 705 301 706
rect 302 705 303 706
rect 303 705 304 706
rect 305 705 306 706
rect 380 580 381 581
rect 382 580 383 581
rect 383 580 384 581
rect 385 580 386 581
rect 380 581 386 585
rect 380 585 381 586
rect 382 585 383 586
rect 383 585 384 586
rect 385 585 386 586
rect 560 1000 561 1001
rect 562 1000 563 1001
rect 563 1000 564 1001
rect 565 1000 566 1001
rect 560 1001 566 1005
rect 560 1005 561 1006
rect 562 1005 563 1006
rect 563 1005 564 1006
rect 565 1005 566 1006
rect 660 920 661 921
rect 662 920 663 921
rect 663 920 664 921
rect 665 920 666 921
rect 660 921 666 925
rect 660 925 661 926
rect 662 925 663 926
rect 663 925 664 926
rect 665 925 666 926
rect 740 360 741 361
rect 742 360 743 361
rect 743 360 744 361
rect 745 360 746 361
rect 740 361 746 365
rect 740 365 741 366
rect 742 365 743 366
rect 743 365 744 366
rect 745 365 746 366
rect 540 580 541 581
rect 542 580 543 581
rect 543 580 544 581
rect 545 580 546 581
rect 540 581 546 585
rect 540 585 541 586
rect 542 585 543 586
rect 543 585 544 586
rect 545 585 546 586
rect 420 880 421 881
rect 422 880 423 881
rect 423 880 424 881
rect 425 880 426 881
rect 420 881 426 885
rect 420 885 421 886
rect 422 885 423 886
rect 423 885 424 886
rect 425 885 426 886
rect 840 480 841 481
rect 842 480 843 481
rect 843 480 844 481
rect 845 480 846 481
rect 840 481 846 485
rect 840 485 841 486
rect 842 485 843 486
rect 843 485 844 486
rect 845 485 846 486
rect 620 500 621 501
rect 622 500 623 501
rect 623 500 624 501
rect 625 500 626 501
rect 620 501 626 505
rect 620 505 621 506
rect 622 505 623 506
rect 623 505 624 506
rect 625 505 626 506
rect 600 740 601 741
rect 602 740 603 741
rect 603 740 604 741
rect 605 740 606 741
rect 600 741 606 745
rect 600 745 601 746
rect 602 745 603 746
rect 603 745 604 746
rect 605 745 606 746
rect 320 780 321 781
rect 322 780 323 781
rect 323 780 324 781
rect 325 780 326 781
rect 320 781 326 785
rect 320 785 321 786
rect 322 785 323 786
rect 323 785 324 786
rect 325 785 326 786
rect 740 980 741 981
rect 742 980 743 981
rect 743 980 744 981
rect 745 980 746 981
rect 740 981 746 985
rect 740 985 741 986
rect 742 985 743 986
rect 743 985 744 986
rect 745 985 746 986
rect 880 860 881 861
rect 882 860 883 861
rect 883 860 884 861
rect 885 860 886 861
rect 880 861 886 865
rect 880 865 881 866
rect 882 865 883 866
rect 883 865 884 866
rect 885 865 886 866
rect 440 620 441 621
rect 442 620 443 621
rect 443 620 444 621
rect 445 620 446 621
rect 440 621 446 625
rect 440 625 441 626
rect 442 625 443 626
rect 443 625 444 626
rect 445 625 446 626
rect 380 560 381 561
rect 382 560 383 561
rect 383 560 384 561
rect 385 560 386 561
rect 380 561 386 565
rect 380 565 381 566
rect 382 565 383 566
rect 383 565 384 566
rect 385 565 386 566
rect 560 980 561 981
rect 562 980 563 981
rect 563 980 564 981
rect 565 980 566 981
rect 560 981 566 985
rect 560 985 561 986
rect 562 985 563 986
rect 563 985 564 986
rect 565 985 566 986
rect 680 400 681 401
rect 682 400 683 401
rect 683 400 684 401
rect 685 400 686 401
rect 680 401 686 405
rect 680 405 681 406
rect 682 405 683 406
rect 683 405 684 406
rect 685 405 686 406
rect 560 400 561 401
rect 562 400 563 401
rect 563 400 564 401
rect 565 400 566 401
rect 560 401 566 405
rect 560 405 561 406
rect 562 405 563 406
rect 563 405 564 406
rect 565 405 566 406
rect 620 780 621 781
rect 622 780 623 781
rect 623 780 624 781
rect 625 780 626 781
rect 620 781 626 785
rect 620 785 621 786
rect 622 785 623 786
rect 623 785 624 786
rect 625 785 626 786
rect 660 1060 661 1061
rect 662 1060 663 1061
rect 663 1060 664 1061
rect 665 1060 666 1061
rect 660 1061 666 1065
rect 660 1065 661 1066
rect 662 1065 663 1066
rect 663 1065 664 1066
rect 665 1065 666 1066
rect 860 640 861 641
rect 862 640 863 641
rect 863 640 864 641
rect 865 640 866 641
rect 860 641 866 645
rect 860 645 861 646
rect 862 645 863 646
rect 863 645 864 646
rect 865 645 866 646
rect 660 640 661 641
rect 662 640 663 641
rect 663 640 664 641
rect 665 640 666 641
rect 660 641 666 645
rect 660 645 661 646
rect 662 645 663 646
rect 663 645 664 646
rect 665 645 666 646
rect 580 380 581 381
rect 582 380 583 381
rect 583 380 584 381
rect 585 380 586 381
rect 580 381 586 385
rect 580 385 581 386
rect 582 385 583 386
rect 583 385 584 386
rect 585 385 586 386
rect 600 460 601 461
rect 602 460 603 461
rect 603 460 604 461
rect 605 460 606 461
rect 600 461 606 465
rect 600 465 601 466
rect 602 465 603 466
rect 603 465 604 466
rect 605 465 606 466
rect 340 660 341 661
rect 342 660 343 661
rect 343 660 344 661
rect 345 660 346 661
rect 340 661 346 665
rect 340 665 341 666
rect 342 665 343 666
rect 343 665 344 666
rect 345 665 346 666
rect 720 1040 721 1041
rect 722 1040 723 1041
rect 723 1040 724 1041
rect 725 1040 726 1041
rect 720 1041 726 1045
rect 720 1045 721 1046
rect 722 1045 723 1046
rect 723 1045 724 1046
rect 725 1045 726 1046
rect 1040 620 1041 621
rect 1042 620 1043 621
rect 1043 620 1044 621
rect 1045 620 1046 621
rect 1040 621 1046 625
rect 1040 625 1041 626
rect 1042 625 1043 626
rect 1043 625 1044 626
rect 1045 625 1046 626
rect 820 840 821 841
rect 822 840 823 841
rect 823 840 824 841
rect 825 840 826 841
rect 820 841 826 845
rect 820 845 821 846
rect 822 845 823 846
rect 823 845 824 846
rect 825 845 826 846
rect 560 840 561 841
rect 562 840 563 841
rect 563 840 564 841
rect 565 840 566 841
rect 560 841 566 845
rect 560 845 561 846
rect 562 845 563 846
rect 563 845 564 846
rect 565 845 566 846
rect 560 460 561 461
rect 562 460 563 461
rect 563 460 564 461
rect 565 460 566 461
rect 560 461 566 465
rect 560 465 561 466
rect 562 465 563 466
rect 563 465 564 466
rect 565 465 566 466
rect 900 860 901 861
rect 902 860 903 861
rect 903 860 904 861
rect 905 860 906 861
rect 900 861 906 865
rect 900 865 901 866
rect 902 865 903 866
rect 903 865 904 866
rect 905 865 906 866
rect 720 440 721 441
rect 722 440 723 441
rect 723 440 724 441
rect 725 440 726 441
rect 720 441 726 445
rect 720 445 721 446
rect 722 445 723 446
rect 723 445 724 446
rect 725 445 726 446
rect 740 880 741 881
rect 742 880 743 881
rect 743 880 744 881
rect 745 880 746 881
rect 740 881 746 885
rect 740 885 741 886
rect 742 885 743 886
rect 743 885 744 886
rect 745 885 746 886
rect 700 400 701 401
rect 702 400 703 401
rect 703 400 704 401
rect 705 400 706 401
rect 700 401 706 405
rect 700 405 701 406
rect 702 405 703 406
rect 703 405 704 406
rect 705 405 706 406
rect 760 1000 761 1001
rect 762 1000 763 1001
rect 763 1000 764 1001
rect 765 1000 766 1001
rect 760 1001 766 1005
rect 760 1005 761 1006
rect 762 1005 763 1006
rect 763 1005 764 1006
rect 765 1005 766 1006
rect 700 460 701 461
rect 702 460 703 461
rect 703 460 704 461
rect 705 460 706 461
rect 700 461 706 465
rect 700 465 701 466
rect 702 465 703 466
rect 703 465 704 466
rect 705 465 706 466
rect 480 400 481 401
rect 482 400 483 401
rect 483 400 484 401
rect 485 400 486 401
rect 480 401 486 405
rect 480 405 481 406
rect 482 405 483 406
rect 483 405 484 406
rect 485 405 486 406
rect 740 560 741 561
rect 742 560 743 561
rect 743 560 744 561
rect 745 560 746 561
rect 740 561 746 565
rect 740 565 741 566
rect 742 565 743 566
rect 743 565 744 566
rect 745 565 746 566
rect 520 860 521 861
rect 522 860 523 861
rect 523 860 524 861
rect 525 860 526 861
rect 520 861 526 865
rect 520 865 521 866
rect 522 865 523 866
rect 523 865 524 866
rect 525 865 526 866
rect 900 540 901 541
rect 902 540 903 541
rect 903 540 904 541
rect 905 540 906 541
rect 900 541 906 545
rect 900 545 901 546
rect 902 545 903 546
rect 903 545 904 546
rect 905 545 906 546
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
<< polysilicon >>
rect 681 699 682 701
rect 684 699 685 701
rect 681 705 682 707
rect 684 705 685 707
rect 581 419 582 421
rect 584 419 585 421
rect 581 425 582 427
rect 584 425 585 427
rect 741 599 742 601
rect 744 599 745 601
rect 741 605 742 607
rect 744 605 745 607
rect 761 519 762 521
rect 764 519 765 521
rect 761 525 762 527
rect 764 525 765 527
rect 641 839 642 841
rect 644 839 645 841
rect 641 845 642 847
rect 644 845 645 847
rect 641 739 642 741
rect 644 739 645 741
rect 641 745 642 747
rect 644 745 645 747
rect 601 919 602 921
rect 604 919 605 921
rect 601 925 602 927
rect 604 925 605 927
rect 501 799 502 801
rect 504 799 505 801
rect 501 805 502 807
rect 504 805 505 807
rect 801 659 802 661
rect 804 659 805 661
rect 801 665 802 667
rect 804 665 805 667
rect 481 639 482 641
rect 484 639 485 641
rect 481 645 482 647
rect 484 645 485 647
rect 841 619 842 621
rect 844 619 845 621
rect 841 625 842 627
rect 844 625 845 627
rect 761 659 762 661
rect 764 659 765 661
rect 761 665 762 667
rect 764 665 765 667
rect 701 699 702 701
rect 704 699 705 701
rect 701 705 702 707
rect 704 705 705 707
rect 521 539 522 541
rect 524 539 525 541
rect 521 545 522 547
rect 524 545 525 547
rect 421 859 422 861
rect 424 859 425 861
rect 421 865 422 867
rect 424 865 425 867
rect 601 899 602 901
rect 604 899 605 901
rect 601 905 602 907
rect 604 905 605 907
rect 441 839 442 841
rect 444 839 445 841
rect 441 845 442 847
rect 444 845 445 847
rect 681 739 682 741
rect 684 739 685 741
rect 681 745 682 747
rect 684 745 685 747
rect 541 539 542 541
rect 544 539 545 541
rect 541 545 542 547
rect 544 545 545 547
rect 861 739 862 741
rect 864 739 865 741
rect 861 745 862 747
rect 864 745 865 747
rect 561 879 562 881
rect 564 879 565 881
rect 561 885 562 887
rect 564 885 565 887
rect 561 599 562 601
rect 564 599 565 601
rect 561 605 562 607
rect 564 605 565 607
rect 641 539 642 541
rect 644 539 645 541
rect 641 545 642 547
rect 644 545 645 547
rect 641 799 642 801
rect 644 799 645 801
rect 641 805 642 807
rect 644 805 645 807
rect 541 799 542 801
rect 544 799 545 801
rect 541 805 542 807
rect 544 805 545 807
rect 581 899 582 901
rect 584 899 585 901
rect 581 905 582 907
rect 584 905 585 907
rect 921 719 922 721
rect 924 719 925 721
rect 921 725 922 727
rect 924 725 925 727
rect 481 759 482 761
rect 484 759 485 761
rect 481 765 482 767
rect 484 765 485 767
rect 681 659 682 661
rect 684 659 685 661
rect 681 665 682 667
rect 684 665 685 667
rect 681 839 682 841
rect 684 839 685 841
rect 681 845 682 847
rect 684 845 685 847
rect 761 479 762 481
rect 764 479 765 481
rect 761 485 762 487
rect 764 485 765 487
rect 401 839 402 841
rect 404 839 405 841
rect 401 845 402 847
rect 404 845 405 847
rect 461 559 462 561
rect 464 559 465 561
rect 461 565 462 567
rect 464 565 465 567
rect 441 719 442 721
rect 444 719 445 721
rect 441 725 442 727
rect 444 725 445 727
rect 601 579 602 581
rect 604 579 605 581
rect 601 585 602 587
rect 604 585 605 587
rect 921 699 922 701
rect 924 699 925 701
rect 921 705 922 707
rect 924 705 925 707
rect 761 619 762 621
rect 764 619 765 621
rect 761 625 762 627
rect 764 625 765 627
rect 701 779 702 781
rect 704 779 705 781
rect 701 785 702 787
rect 704 785 705 787
rect 641 639 642 641
rect 644 639 645 641
rect 641 645 642 647
rect 644 645 645 647
rect 441 699 442 701
rect 444 699 445 701
rect 441 705 442 707
rect 444 705 445 707
rect 601 639 602 641
rect 604 639 605 641
rect 601 645 602 647
rect 604 645 605 647
rect 721 599 722 601
rect 724 599 725 601
rect 721 605 722 607
rect 724 605 725 607
rect 441 899 442 901
rect 444 899 445 901
rect 441 905 442 907
rect 444 905 445 907
rect 601 519 602 521
rect 604 519 605 521
rect 601 525 602 527
rect 604 525 605 527
rect 581 679 582 681
rect 584 679 585 681
rect 581 685 582 687
rect 584 685 585 687
rect 721 679 722 681
rect 724 679 725 681
rect 721 685 722 687
rect 724 685 725 687
rect 801 699 802 701
rect 804 699 805 701
rect 801 705 802 707
rect 804 705 805 707
rect 781 579 782 581
rect 784 579 785 581
rect 781 585 782 587
rect 784 585 785 587
rect 861 599 862 601
rect 864 599 865 601
rect 861 605 862 607
rect 864 605 865 607
rect 501 939 502 941
rect 504 939 505 941
rect 501 945 502 947
rect 504 945 505 947
rect 741 719 742 721
rect 744 719 745 721
rect 741 725 742 727
rect 744 725 745 727
rect 521 759 522 761
rect 524 759 525 761
rect 521 765 522 767
rect 524 765 525 767
rect 841 739 842 741
rect 844 739 845 741
rect 841 745 842 747
rect 844 745 845 747
rect 701 579 702 581
rect 704 579 705 581
rect 701 585 702 587
rect 704 585 705 587
rect 581 539 582 541
rect 584 539 585 541
rect 581 545 582 547
rect 584 545 585 547
rect 781 759 782 761
rect 784 759 785 761
rect 781 765 782 767
rect 784 765 785 767
rect 601 839 602 841
rect 604 839 605 841
rect 601 845 602 847
rect 604 845 605 847
rect 661 439 662 441
rect 664 439 665 441
rect 661 445 662 447
rect 664 445 665 447
rect 781 639 782 641
rect 784 639 785 641
rect 781 645 782 647
rect 784 645 785 647
rect 521 679 522 681
rect 524 679 525 681
rect 521 685 522 687
rect 524 685 525 687
rect 341 679 342 681
rect 344 679 345 681
rect 341 685 342 687
rect 344 685 345 687
rect 481 659 482 661
rect 484 659 485 661
rect 481 665 482 667
rect 484 665 485 667
rect 601 979 602 981
rect 604 979 605 981
rect 601 985 602 987
rect 604 985 605 987
rect 681 599 682 601
rect 684 599 685 601
rect 681 605 682 607
rect 684 605 685 607
rect 681 899 682 901
rect 684 899 685 901
rect 681 905 682 907
rect 684 905 685 907
rect 821 899 822 901
rect 824 899 825 901
rect 821 905 822 907
rect 824 905 825 907
rect 661 779 662 781
rect 664 779 665 781
rect 661 785 662 787
rect 664 785 665 787
rect 681 859 682 861
rect 684 859 685 861
rect 681 865 682 867
rect 684 865 685 867
rect 661 879 662 881
rect 664 879 665 881
rect 661 885 662 887
rect 664 885 665 887
rect 341 699 342 701
rect 344 699 345 701
rect 341 705 342 707
rect 344 705 345 707
rect 541 559 542 561
rect 544 559 545 561
rect 541 565 542 567
rect 544 565 545 567
rect 381 859 382 861
rect 384 859 385 861
rect 381 865 382 867
rect 384 865 385 867
rect 721 739 722 741
rect 724 739 725 741
rect 721 745 722 747
rect 724 745 725 747
rect 521 739 522 741
rect 524 739 525 741
rect 521 745 522 747
rect 524 745 525 747
rect 621 879 622 881
rect 624 879 625 881
rect 621 885 622 887
rect 624 885 625 887
rect 621 379 622 381
rect 624 379 625 381
rect 621 385 622 387
rect 624 385 625 387
rect 661 619 662 621
rect 664 619 665 621
rect 661 625 662 627
rect 664 625 665 627
rect 761 699 762 701
rect 764 699 765 701
rect 761 705 762 707
rect 764 705 765 707
rect 861 499 862 501
rect 864 499 865 501
rect 861 505 862 507
rect 864 505 865 507
rect 501 839 502 841
rect 504 839 505 841
rect 501 845 502 847
rect 504 845 505 847
rect 701 479 702 481
rect 704 479 705 481
rect 701 485 702 487
rect 704 485 705 487
rect 521 559 522 561
rect 524 559 525 561
rect 521 565 522 567
rect 524 565 525 567
rect 961 679 962 681
rect 964 679 965 681
rect 961 685 962 687
rect 964 685 965 687
rect 441 559 442 561
rect 444 559 445 561
rect 441 565 442 567
rect 444 565 445 567
rect 481 779 482 781
rect 484 779 485 781
rect 481 785 482 787
rect 484 785 485 787
rect 481 879 482 881
rect 484 879 485 881
rect 481 885 482 887
rect 484 885 485 887
rect 661 679 662 681
rect 664 679 665 681
rect 661 685 662 687
rect 664 685 665 687
rect 641 459 642 461
rect 644 459 645 461
rect 641 465 642 467
rect 644 465 645 467
rect 841 839 842 841
rect 844 839 845 841
rect 841 845 842 847
rect 844 845 845 847
rect 621 679 622 681
rect 624 679 625 681
rect 621 685 622 687
rect 624 685 625 687
rect 921 779 922 781
rect 924 779 925 781
rect 921 785 922 787
rect 924 785 925 787
rect 441 639 442 641
rect 444 639 445 641
rect 441 645 442 647
rect 444 645 445 647
rect 921 799 922 801
rect 924 799 925 801
rect 921 805 922 807
rect 924 805 925 807
rect 381 599 382 601
rect 384 599 385 601
rect 381 605 382 607
rect 384 605 385 607
rect 801 819 802 821
rect 804 819 805 821
rect 801 825 802 827
rect 804 825 805 827
rect 461 919 462 921
rect 464 919 465 921
rect 461 925 462 927
rect 464 925 465 927
rect 361 539 362 541
rect 364 539 365 541
rect 361 545 362 547
rect 364 545 365 547
rect 661 559 662 561
rect 664 559 665 561
rect 661 565 662 567
rect 664 565 665 567
rect 641 479 642 481
rect 644 479 645 481
rect 641 485 642 487
rect 644 485 645 487
rect 741 619 742 621
rect 744 619 745 621
rect 741 625 742 627
rect 744 625 745 627
rect 661 899 662 901
rect 664 899 665 901
rect 661 905 662 907
rect 664 905 665 907
rect 801 479 802 481
rect 804 479 805 481
rect 801 485 802 487
rect 804 485 805 487
rect 801 719 802 721
rect 804 719 805 721
rect 801 725 802 727
rect 804 725 805 727
rect 461 619 462 621
rect 464 619 465 621
rect 461 625 462 627
rect 464 625 465 627
rect 561 539 562 541
rect 564 539 565 541
rect 561 545 562 547
rect 564 545 565 547
rect 621 719 622 721
rect 624 719 625 721
rect 621 725 622 727
rect 624 725 625 727
rect 801 799 802 801
rect 804 799 805 801
rect 801 805 802 807
rect 804 805 805 807
rect 601 599 602 601
rect 604 599 605 601
rect 601 605 602 607
rect 604 605 605 607
rect 921 839 922 841
rect 924 839 925 841
rect 921 845 922 847
rect 924 845 925 847
rect 481 539 482 541
rect 484 539 485 541
rect 481 545 482 547
rect 484 545 485 547
rect 921 559 922 561
rect 924 559 925 561
rect 921 565 922 567
rect 924 565 925 567
rect 641 699 642 701
rect 644 699 645 701
rect 641 705 642 707
rect 644 705 645 707
rect 641 519 642 521
rect 644 519 645 521
rect 641 525 642 527
rect 644 525 645 527
rect 921 679 922 681
rect 924 679 925 681
rect 921 685 922 687
rect 924 685 925 687
rect 621 759 622 761
rect 624 759 625 761
rect 621 765 622 767
rect 624 765 625 767
rect 421 739 422 741
rect 424 739 425 741
rect 421 745 422 747
rect 424 745 425 747
rect 801 519 802 521
rect 804 519 805 521
rect 801 525 802 527
rect 804 525 805 527
rect 721 459 722 461
rect 724 459 725 461
rect 721 465 722 467
rect 724 465 725 467
rect 921 579 922 581
rect 924 579 925 581
rect 921 585 922 587
rect 924 585 925 587
rect 561 779 562 781
rect 564 779 565 781
rect 561 785 562 787
rect 564 785 565 787
rect 501 379 502 381
rect 504 379 505 381
rect 501 385 502 387
rect 504 385 505 387
rect 941 599 942 601
rect 944 599 945 601
rect 941 605 942 607
rect 944 605 945 607
rect 421 539 422 541
rect 424 539 425 541
rect 421 545 422 547
rect 424 545 425 547
rect 941 619 942 621
rect 944 619 945 621
rect 941 625 942 627
rect 944 625 945 627
rect 561 719 562 721
rect 564 719 565 721
rect 561 725 562 727
rect 564 725 565 727
rect 461 859 462 861
rect 464 859 465 861
rect 461 865 462 867
rect 464 865 465 867
rect 561 819 562 821
rect 564 819 565 821
rect 561 825 562 827
rect 564 825 565 827
rect 741 639 742 641
rect 744 639 745 641
rect 741 645 742 647
rect 744 645 745 647
rect 761 879 762 881
rect 764 879 765 881
rect 761 885 762 887
rect 764 885 765 887
rect 481 679 482 681
rect 484 679 485 681
rect 481 685 482 687
rect 484 685 485 687
rect 841 939 842 941
rect 844 939 845 941
rect 841 945 842 947
rect 844 945 845 947
rect 861 459 862 461
rect 864 459 865 461
rect 861 465 862 467
rect 864 465 865 467
rect 661 599 662 601
rect 664 599 665 601
rect 661 605 662 607
rect 664 605 665 607
rect 481 479 482 481
rect 484 479 485 481
rect 481 485 482 487
rect 484 485 485 487
rect 721 519 722 521
rect 724 519 725 521
rect 721 525 722 527
rect 724 525 725 527
rect 501 579 502 581
rect 504 579 505 581
rect 501 585 502 587
rect 504 585 505 587
rect 361 839 362 841
rect 364 839 365 841
rect 361 845 362 847
rect 364 845 365 847
rect 361 819 362 821
rect 364 819 365 821
rect 361 825 362 827
rect 364 825 365 827
rect 741 519 742 521
rect 744 519 745 521
rect 741 525 742 527
rect 744 525 745 527
rect 841 779 842 781
rect 844 779 845 781
rect 841 785 842 787
rect 844 785 845 787
rect 381 619 382 621
rect 384 619 385 621
rect 381 625 382 627
rect 384 625 385 627
rect 481 839 482 841
rect 484 839 485 841
rect 481 845 482 847
rect 484 845 485 847
rect 561 479 562 481
rect 564 479 565 481
rect 561 485 562 487
rect 564 485 565 487
rect 441 679 442 681
rect 444 679 445 681
rect 441 685 442 687
rect 444 685 445 687
rect 501 699 502 701
rect 504 699 505 701
rect 501 705 502 707
rect 504 705 505 707
rect 521 839 522 841
rect 524 839 525 841
rect 521 845 522 847
rect 524 845 525 847
rect 541 639 542 641
rect 544 639 545 641
rect 541 645 542 647
rect 544 645 545 647
rect 801 559 802 561
rect 804 559 805 561
rect 801 565 802 567
rect 804 565 805 567
rect 561 519 562 521
rect 564 519 565 521
rect 561 525 562 527
rect 564 525 565 527
rect 581 699 582 701
rect 584 699 585 701
rect 581 705 582 707
rect 584 705 585 707
rect 601 799 602 801
rect 604 799 605 801
rect 601 805 602 807
rect 604 805 605 807
rect 821 879 822 881
rect 824 879 825 881
rect 821 885 822 887
rect 824 885 825 887
rect 761 779 762 781
rect 764 779 765 781
rect 761 785 762 787
rect 764 785 765 787
rect 621 959 622 961
rect 624 959 625 961
rect 621 965 622 967
rect 624 965 625 967
rect 481 699 482 701
rect 484 699 485 701
rect 481 705 482 707
rect 484 705 485 707
rect 501 439 502 441
rect 504 439 505 441
rect 501 445 502 447
rect 504 445 505 447
rect 521 639 522 641
rect 524 639 525 641
rect 521 645 522 647
rect 524 645 525 647
rect 761 679 762 681
rect 764 679 765 681
rect 761 685 762 687
rect 764 685 765 687
rect 541 819 542 821
rect 544 819 545 821
rect 541 825 542 827
rect 544 825 545 827
rect 561 379 562 381
rect 564 379 565 381
rect 561 385 562 387
rect 564 385 565 387
rect 861 779 862 781
rect 864 779 865 781
rect 861 785 862 787
rect 864 785 865 787
rect 661 459 662 461
rect 664 459 665 461
rect 661 465 662 467
rect 664 465 665 467
rect 681 299 682 301
rect 684 299 685 301
rect 681 305 682 307
rect 684 305 685 307
rect 641 619 642 621
rect 644 619 645 621
rect 641 625 642 627
rect 644 625 645 627
rect 561 659 562 661
rect 564 659 565 661
rect 561 665 562 667
rect 564 665 565 667
rect 361 599 362 601
rect 364 599 365 601
rect 361 605 362 607
rect 364 605 365 607
rect 641 1019 642 1021
rect 644 1019 645 1021
rect 641 1025 642 1027
rect 644 1025 645 1027
rect 721 819 722 821
rect 724 819 725 821
rect 721 825 722 827
rect 724 825 725 827
rect 761 719 762 721
rect 764 719 765 721
rect 761 725 762 727
rect 764 725 765 727
rect 661 799 662 801
rect 664 799 665 801
rect 661 805 662 807
rect 664 805 665 807
rect 561 679 562 681
rect 564 679 565 681
rect 561 685 562 687
rect 564 685 565 687
rect 461 739 462 741
rect 464 739 465 741
rect 461 745 462 747
rect 464 745 465 747
rect 741 319 742 321
rect 744 319 745 321
rect 741 325 742 327
rect 744 325 745 327
rect 701 519 702 521
rect 704 519 705 521
rect 701 525 702 527
rect 704 525 705 527
rect 501 719 502 721
rect 504 719 505 721
rect 501 725 502 727
rect 504 725 505 727
rect 701 899 702 901
rect 704 899 705 901
rect 701 905 702 907
rect 704 905 705 907
rect 961 579 962 581
rect 964 579 965 581
rect 961 585 962 587
rect 964 585 965 587
rect 741 959 742 961
rect 744 959 745 961
rect 741 965 742 967
rect 744 965 745 967
rect 601 1039 602 1041
rect 604 1039 605 1041
rect 601 1045 602 1047
rect 604 1045 605 1047
rect 761 939 762 941
rect 764 939 765 941
rect 761 945 762 947
rect 764 945 765 947
rect 801 639 802 641
rect 804 639 805 641
rect 801 645 802 647
rect 804 645 805 647
rect 321 759 322 761
rect 324 759 325 761
rect 321 765 322 767
rect 324 765 325 767
rect 821 599 822 601
rect 824 599 825 601
rect 821 605 822 607
rect 824 605 825 607
rect 721 299 722 301
rect 724 299 725 301
rect 721 305 722 307
rect 724 305 725 307
rect 681 459 682 461
rect 684 459 685 461
rect 681 465 682 467
rect 684 465 685 467
rect 821 559 822 561
rect 824 559 825 561
rect 821 565 822 567
rect 824 565 825 567
rect 721 799 722 801
rect 724 799 725 801
rect 721 805 722 807
rect 724 805 725 807
rect 621 919 622 921
rect 624 919 625 921
rect 621 925 622 927
rect 624 925 625 927
rect 361 799 362 801
rect 364 799 365 801
rect 361 805 362 807
rect 364 805 365 807
rect 541 759 542 761
rect 544 759 545 761
rect 541 765 542 767
rect 544 765 545 767
rect 481 499 482 501
rect 484 499 485 501
rect 481 505 482 507
rect 484 505 485 507
rect 621 559 622 561
rect 624 559 625 561
rect 621 565 622 567
rect 624 565 625 567
rect 701 1019 702 1021
rect 704 1019 705 1021
rect 701 1025 702 1027
rect 704 1025 705 1027
rect 861 919 862 921
rect 864 919 865 921
rect 861 925 862 927
rect 864 925 865 927
rect 861 759 862 761
rect 864 759 865 761
rect 861 765 862 767
rect 864 765 865 767
rect 981 679 982 681
rect 984 679 985 681
rect 981 685 982 687
rect 984 685 985 687
rect 421 839 422 841
rect 424 839 425 841
rect 421 845 422 847
rect 424 845 425 847
rect 781 839 782 841
rect 784 839 785 841
rect 781 845 782 847
rect 784 845 785 847
rect 841 459 842 461
rect 844 459 845 461
rect 841 465 842 467
rect 844 465 845 467
rect 501 779 502 781
rect 504 779 505 781
rect 501 785 502 787
rect 504 785 505 787
rect 581 599 582 601
rect 584 599 585 601
rect 581 605 582 607
rect 584 605 585 607
rect 701 319 702 321
rect 704 319 705 321
rect 701 325 702 327
rect 704 325 705 327
rect 561 359 562 361
rect 564 359 565 361
rect 561 365 562 367
rect 564 365 565 367
rect 781 899 782 901
rect 784 899 785 901
rect 781 905 782 907
rect 784 905 785 907
rect 481 439 482 441
rect 484 439 485 441
rect 481 445 482 447
rect 484 445 485 447
rect 801 539 802 541
rect 804 539 805 541
rect 801 545 802 547
rect 804 545 805 547
rect 761 359 762 361
rect 764 359 765 361
rect 761 365 762 367
rect 764 365 765 367
rect 621 479 622 481
rect 624 479 625 481
rect 621 485 622 487
rect 624 485 625 487
rect 841 679 842 681
rect 844 679 845 681
rect 841 685 842 687
rect 844 685 845 687
rect 561 739 562 741
rect 564 739 565 741
rect 561 745 562 747
rect 564 745 565 747
rect 901 619 902 621
rect 904 619 905 621
rect 901 625 902 627
rect 904 625 905 627
rect 441 479 442 481
rect 444 479 445 481
rect 441 485 442 487
rect 444 485 445 487
rect 761 399 762 401
rect 764 399 765 401
rect 761 405 762 407
rect 764 405 765 407
rect 541 719 542 721
rect 544 719 545 721
rect 541 725 542 727
rect 544 725 545 727
rect 661 819 662 821
rect 664 819 665 821
rect 661 825 662 827
rect 664 825 665 827
rect 401 639 402 641
rect 404 639 405 641
rect 401 645 402 647
rect 404 645 405 647
rect 741 1019 742 1021
rect 744 1019 745 1021
rect 741 1025 742 1027
rect 744 1025 745 1027
rect 541 999 542 1001
rect 544 999 545 1001
rect 541 1005 542 1007
rect 544 1005 545 1007
rect 781 399 782 401
rect 784 399 785 401
rect 781 405 782 407
rect 784 405 785 407
rect 661 1039 662 1041
rect 664 1039 665 1041
rect 661 1045 662 1047
rect 664 1045 665 1047
rect 601 1059 602 1061
rect 604 1059 605 1061
rect 601 1065 602 1067
rect 604 1065 605 1067
rect 481 739 482 741
rect 484 739 485 741
rect 481 745 482 747
rect 484 745 485 747
rect 461 639 462 641
rect 464 639 465 641
rect 461 645 462 647
rect 464 645 465 647
rect 461 899 462 901
rect 464 899 465 901
rect 461 905 462 907
rect 464 905 465 907
rect 581 459 582 461
rect 584 459 585 461
rect 581 465 582 467
rect 584 465 585 467
rect 641 399 642 401
rect 644 399 645 401
rect 641 405 642 407
rect 644 405 645 407
rect 961 759 962 761
rect 964 759 965 761
rect 961 765 962 767
rect 964 765 965 767
rect 561 959 562 961
rect 564 959 565 961
rect 561 965 562 967
rect 564 965 565 967
rect 681 259 682 261
rect 684 259 685 261
rect 681 265 682 267
rect 684 265 685 267
rect 561 579 562 581
rect 564 579 565 581
rect 561 585 562 587
rect 564 585 565 587
rect 681 919 682 921
rect 684 919 685 921
rect 681 925 682 927
rect 684 925 685 927
rect 501 959 502 961
rect 504 959 505 961
rect 501 965 502 967
rect 504 965 505 967
rect 621 319 622 321
rect 624 319 625 321
rect 621 325 622 327
rect 624 325 625 327
rect 601 379 602 381
rect 604 379 605 381
rect 601 385 602 387
rect 604 385 605 387
rect 881 479 882 481
rect 884 479 885 481
rect 881 485 882 487
rect 884 485 885 487
rect 1001 779 1002 781
rect 1004 779 1005 781
rect 1001 785 1002 787
rect 1004 785 1005 787
rect 261 719 262 721
rect 264 719 265 721
rect 261 725 262 727
rect 264 725 265 727
rect 561 419 562 421
rect 564 419 565 421
rect 561 425 562 427
rect 564 425 565 427
rect 261 739 262 741
rect 264 739 265 741
rect 261 745 262 747
rect 264 745 265 747
rect 861 839 862 841
rect 864 839 865 841
rect 861 845 862 847
rect 864 845 865 847
rect 461 719 462 721
rect 464 719 465 721
rect 461 725 462 727
rect 464 725 465 727
rect 641 719 642 721
rect 644 719 645 721
rect 641 725 642 727
rect 644 725 645 727
rect 721 359 722 361
rect 724 359 725 361
rect 721 365 722 367
rect 724 365 725 367
rect 801 459 802 461
rect 804 459 805 461
rect 801 465 802 467
rect 804 465 805 467
rect 781 879 782 881
rect 784 879 785 881
rect 781 885 782 887
rect 784 885 785 887
rect 901 879 902 881
rect 904 879 905 881
rect 901 885 902 887
rect 904 885 905 887
rect 781 459 782 461
rect 784 459 785 461
rect 781 465 782 467
rect 784 465 785 467
rect 621 1039 622 1041
rect 624 1039 625 1041
rect 621 1045 622 1047
rect 624 1045 625 1047
rect 681 679 682 681
rect 684 679 685 681
rect 681 685 682 687
rect 684 685 685 687
rect 781 539 782 541
rect 784 539 785 541
rect 781 545 782 547
rect 784 545 785 547
rect 701 959 702 961
rect 704 959 705 961
rect 701 965 702 967
rect 704 965 705 967
rect 621 979 622 981
rect 624 979 625 981
rect 621 985 622 987
rect 624 985 625 987
rect 721 639 722 641
rect 724 639 725 641
rect 721 645 722 647
rect 724 645 725 647
rect 701 739 702 741
rect 704 739 705 741
rect 701 745 702 747
rect 704 745 705 747
rect 581 1019 582 1021
rect 584 1019 585 1021
rect 581 1025 582 1027
rect 584 1025 585 1027
rect 261 639 262 641
rect 264 639 265 641
rect 261 645 262 647
rect 264 645 265 647
rect 501 919 502 921
rect 504 919 505 921
rect 501 925 502 927
rect 504 925 505 927
rect 741 459 742 461
rect 744 459 745 461
rect 741 465 742 467
rect 744 465 745 467
rect 281 739 282 741
rect 284 739 285 741
rect 281 745 282 747
rect 284 745 285 747
rect 341 799 342 801
rect 344 799 345 801
rect 341 805 342 807
rect 344 805 345 807
rect 621 399 622 401
rect 624 399 625 401
rect 621 405 622 407
rect 624 405 625 407
rect 781 439 782 441
rect 784 439 785 441
rect 781 445 782 447
rect 784 445 785 447
rect 361 639 362 641
rect 364 639 365 641
rect 361 645 362 647
rect 364 645 365 647
rect 401 659 402 661
rect 404 659 405 661
rect 401 665 402 667
rect 404 665 405 667
rect 521 919 522 921
rect 524 919 525 921
rect 521 925 522 927
rect 524 925 525 927
rect 721 659 722 661
rect 724 659 725 661
rect 721 665 722 667
rect 724 665 725 667
rect 981 759 982 761
rect 984 759 985 761
rect 981 765 982 767
rect 984 765 985 767
rect 901 839 902 841
rect 904 839 905 841
rect 901 845 902 847
rect 904 845 905 847
rect 601 339 602 341
rect 604 339 605 341
rect 601 345 602 347
rect 604 345 605 347
rect 981 559 982 561
rect 984 559 985 561
rect 981 565 982 567
rect 984 565 985 567
rect 681 639 682 641
rect 684 639 685 641
rect 681 645 682 647
rect 684 645 685 647
rect 361 579 362 581
rect 364 579 365 581
rect 361 585 362 587
rect 364 585 365 587
rect 601 679 602 681
rect 604 679 605 681
rect 601 685 602 687
rect 604 685 605 687
rect 921 859 922 861
rect 924 859 925 861
rect 921 865 922 867
rect 924 865 925 867
rect 321 699 322 701
rect 324 699 325 701
rect 321 705 322 707
rect 324 705 325 707
rect 581 779 582 781
rect 584 779 585 781
rect 581 785 582 787
rect 584 785 585 787
rect 701 679 702 681
rect 704 679 705 681
rect 701 685 702 687
rect 704 685 705 687
rect 721 959 722 961
rect 724 959 725 961
rect 721 965 722 967
rect 724 965 725 967
rect 341 739 342 741
rect 344 739 345 741
rect 341 745 342 747
rect 344 745 345 747
rect 601 479 602 481
rect 604 479 605 481
rect 601 485 602 487
rect 604 485 605 487
rect 561 339 562 341
rect 564 339 565 341
rect 561 345 562 347
rect 564 345 565 347
rect 701 799 702 801
rect 704 799 705 801
rect 701 805 702 807
rect 704 805 705 807
rect 941 579 942 581
rect 944 579 945 581
rect 941 585 942 587
rect 944 585 945 587
rect 481 459 482 461
rect 484 459 485 461
rect 481 465 482 467
rect 484 465 485 467
rect 421 479 422 481
rect 424 479 425 481
rect 421 485 422 487
rect 424 485 425 487
rect 481 519 482 521
rect 484 519 485 521
rect 481 525 482 527
rect 484 525 485 527
rect 641 279 642 281
rect 644 279 645 281
rect 641 285 642 287
rect 644 285 645 287
rect 881 599 882 601
rect 884 599 885 601
rect 881 605 882 607
rect 884 605 885 607
rect 641 819 642 821
rect 644 819 645 821
rect 641 825 642 827
rect 644 825 645 827
rect 721 719 722 721
rect 724 719 725 721
rect 721 725 722 727
rect 724 725 725 727
rect 381 539 382 541
rect 384 539 385 541
rect 381 545 382 547
rect 384 545 385 547
rect 441 599 442 601
rect 444 599 445 601
rect 441 605 442 607
rect 444 605 445 607
rect 761 499 762 501
rect 764 499 765 501
rect 761 505 762 507
rect 764 505 765 507
rect 601 419 602 421
rect 604 419 605 421
rect 601 425 602 427
rect 604 425 605 427
rect 621 579 622 581
rect 624 579 625 581
rect 621 585 622 587
rect 624 585 625 587
rect 701 359 702 361
rect 704 359 705 361
rect 701 365 702 367
rect 704 365 705 367
rect 941 539 942 541
rect 944 539 945 541
rect 941 545 942 547
rect 944 545 945 547
rect 341 759 342 761
rect 344 759 345 761
rect 341 765 342 767
rect 344 765 345 767
rect 581 799 582 801
rect 584 799 585 801
rect 581 805 582 807
rect 584 805 585 807
rect 501 659 502 661
rect 504 659 505 661
rect 501 665 502 667
rect 504 665 505 667
rect 501 519 502 521
rect 504 519 505 521
rect 501 525 502 527
rect 504 525 505 527
rect 661 319 662 321
rect 664 319 665 321
rect 661 325 662 327
rect 664 325 665 327
rect 501 599 502 601
rect 504 599 505 601
rect 501 605 502 607
rect 504 605 505 607
rect 661 419 662 421
rect 664 419 665 421
rect 661 425 662 427
rect 664 425 665 427
rect 621 1059 622 1061
rect 624 1059 625 1061
rect 621 1065 622 1067
rect 624 1065 625 1067
rect 521 519 522 521
rect 524 519 525 521
rect 521 525 522 527
rect 524 525 525 527
rect 481 799 482 801
rect 484 799 485 801
rect 481 805 482 807
rect 484 805 485 807
rect 461 539 462 541
rect 464 539 465 541
rect 461 545 462 547
rect 464 545 465 547
rect 721 939 722 941
rect 724 939 725 941
rect 721 945 722 947
rect 724 945 725 947
rect 901 579 902 581
rect 904 579 905 581
rect 901 585 902 587
rect 904 585 905 587
rect 301 659 302 661
rect 304 659 305 661
rect 301 665 302 667
rect 304 665 305 667
rect 521 419 522 421
rect 524 419 525 421
rect 521 425 522 427
rect 524 425 525 427
rect 681 979 682 981
rect 684 979 685 981
rect 681 985 682 987
rect 684 985 685 987
rect 421 679 422 681
rect 424 679 425 681
rect 421 685 422 687
rect 424 685 425 687
rect 621 839 622 841
rect 624 839 625 841
rect 621 845 622 847
rect 624 845 625 847
rect 981 699 982 701
rect 984 699 985 701
rect 981 705 982 707
rect 984 705 985 707
rect 321 619 322 621
rect 324 619 325 621
rect 321 625 322 627
rect 324 625 325 627
rect 381 639 382 641
rect 384 639 385 641
rect 381 645 382 647
rect 384 645 385 647
rect 741 539 742 541
rect 744 539 745 541
rect 741 545 742 547
rect 744 545 745 547
rect 401 619 402 621
rect 404 619 405 621
rect 401 625 402 627
rect 404 625 405 627
rect 581 639 582 641
rect 584 639 585 641
rect 581 645 582 647
rect 584 645 585 647
rect 621 1019 622 1021
rect 624 1019 625 1021
rect 621 1025 622 1027
rect 624 1025 625 1027
rect 721 479 722 481
rect 724 479 725 481
rect 721 485 722 487
rect 724 485 725 487
rect 341 579 342 581
rect 344 579 345 581
rect 341 585 342 587
rect 344 585 345 587
rect 881 639 882 641
rect 884 639 885 641
rect 881 645 882 647
rect 884 645 885 647
rect 581 399 582 401
rect 584 399 585 401
rect 581 405 582 407
rect 584 405 585 407
rect 821 699 822 701
rect 824 699 825 701
rect 821 705 822 707
rect 824 705 825 707
rect 501 759 502 761
rect 504 759 505 761
rect 501 765 502 767
rect 504 765 505 767
rect 441 879 442 881
rect 444 879 445 881
rect 441 885 442 887
rect 444 885 445 887
rect 761 439 762 441
rect 764 439 765 441
rect 761 445 762 447
rect 764 445 765 447
rect 601 299 602 301
rect 604 299 605 301
rect 601 305 602 307
rect 604 305 605 307
rect 961 699 962 701
rect 964 699 965 701
rect 961 705 962 707
rect 964 705 965 707
rect 541 699 542 701
rect 544 699 545 701
rect 541 705 542 707
rect 544 705 545 707
rect 841 899 842 901
rect 844 899 845 901
rect 841 905 842 907
rect 844 905 845 907
rect 561 859 562 861
rect 564 859 565 861
rect 561 865 562 867
rect 564 865 565 867
rect 681 439 682 441
rect 684 439 685 441
rect 681 445 682 447
rect 684 445 685 447
rect 801 879 802 881
rect 804 879 805 881
rect 801 885 802 887
rect 804 885 805 887
rect 781 519 782 521
rect 784 519 785 521
rect 781 525 782 527
rect 784 525 785 527
rect 401 759 402 761
rect 404 759 405 761
rect 401 765 402 767
rect 404 765 405 767
rect 721 279 722 281
rect 724 279 725 281
rect 721 285 722 287
rect 724 285 725 287
rect 501 619 502 621
rect 504 619 505 621
rect 501 625 502 627
rect 504 625 505 627
rect 461 499 462 501
rect 464 499 465 501
rect 461 505 462 507
rect 464 505 465 507
rect 841 719 842 721
rect 844 719 845 721
rect 841 725 842 727
rect 844 725 845 727
rect 621 999 622 1001
rect 624 999 625 1001
rect 621 1005 622 1007
rect 624 1005 625 1007
rect 661 999 662 1001
rect 664 999 665 1001
rect 661 1005 662 1007
rect 664 1005 665 1007
rect 561 639 562 641
rect 564 639 565 641
rect 561 645 562 647
rect 564 645 565 647
rect 261 599 262 601
rect 264 599 265 601
rect 261 605 262 607
rect 264 605 265 607
rect 401 559 402 561
rect 404 559 405 561
rect 401 565 402 567
rect 404 565 405 567
rect 421 659 422 661
rect 424 659 425 661
rect 421 665 422 667
rect 424 665 425 667
rect 261 659 262 661
rect 264 659 265 661
rect 261 665 262 667
rect 264 665 265 667
rect 661 759 662 761
rect 664 759 665 761
rect 661 765 662 767
rect 664 765 665 767
rect 1021 639 1022 641
rect 1024 639 1025 641
rect 1021 645 1022 647
rect 1024 645 1025 647
rect 641 959 642 961
rect 644 959 645 961
rect 641 965 642 967
rect 644 965 645 967
rect 301 759 302 761
rect 304 759 305 761
rect 301 765 302 767
rect 304 765 305 767
rect 661 859 662 861
rect 664 859 665 861
rect 661 865 662 867
rect 664 865 665 867
rect 961 539 962 541
rect 964 539 965 541
rect 961 545 962 547
rect 964 545 965 547
rect 821 779 822 781
rect 824 779 825 781
rect 821 785 822 787
rect 824 785 825 787
rect 841 879 842 881
rect 844 879 845 881
rect 841 885 842 887
rect 844 885 845 887
rect 741 499 742 501
rect 744 499 745 501
rect 741 505 742 507
rect 744 505 745 507
rect 621 419 622 421
rect 624 419 625 421
rect 621 425 622 427
rect 624 425 625 427
rect 881 899 882 901
rect 884 899 885 901
rect 881 905 882 907
rect 884 905 885 907
rect 281 619 282 621
rect 284 619 285 621
rect 281 625 282 627
rect 284 625 285 627
rect 641 339 642 341
rect 644 339 645 341
rect 641 345 642 347
rect 644 345 645 347
rect 541 619 542 621
rect 544 619 545 621
rect 541 625 542 627
rect 544 625 545 627
rect 481 619 482 621
rect 484 619 485 621
rect 481 625 482 627
rect 484 625 485 627
rect 481 419 482 421
rect 484 419 485 421
rect 481 425 482 427
rect 484 425 485 427
rect 241 679 242 681
rect 244 679 245 681
rect 241 685 242 687
rect 244 685 245 687
rect 601 819 602 821
rect 604 819 605 821
rect 601 825 602 827
rect 604 825 605 827
rect 561 619 562 621
rect 564 619 565 621
rect 561 625 562 627
rect 564 625 565 627
rect 901 819 902 821
rect 904 819 905 821
rect 901 825 902 827
rect 904 825 905 827
rect 801 939 802 941
rect 804 939 805 941
rect 801 945 802 947
rect 804 945 805 947
rect 821 479 822 481
rect 824 479 825 481
rect 821 485 822 487
rect 824 485 825 487
rect 1001 699 1002 701
rect 1004 699 1005 701
rect 1001 705 1002 707
rect 1004 705 1005 707
rect 321 679 322 681
rect 324 679 325 681
rect 321 685 322 687
rect 324 685 325 687
rect 741 379 742 381
rect 744 379 745 381
rect 741 385 742 387
rect 744 385 745 387
rect 941 819 942 821
rect 944 819 945 821
rect 941 825 942 827
rect 944 825 945 827
rect 741 1039 742 1041
rect 744 1039 745 1041
rect 741 1045 742 1047
rect 744 1045 745 1047
rect 421 519 422 521
rect 424 519 425 521
rect 421 525 422 527
rect 424 525 425 527
rect 781 939 782 941
rect 784 939 785 941
rect 781 945 782 947
rect 784 945 785 947
rect 901 479 902 481
rect 904 479 905 481
rect 901 485 902 487
rect 904 485 905 487
rect 741 399 742 401
rect 744 399 745 401
rect 741 405 742 407
rect 744 405 745 407
rect 881 759 882 761
rect 884 759 885 761
rect 881 765 882 767
rect 884 765 885 767
rect 701 999 702 1001
rect 704 999 705 1001
rect 701 1005 702 1007
rect 704 1005 705 1007
rect 641 559 642 561
rect 644 559 645 561
rect 641 565 642 567
rect 644 565 645 567
rect 601 319 602 321
rect 604 319 605 321
rect 601 325 602 327
rect 604 325 605 327
rect 761 379 762 381
rect 764 379 765 381
rect 761 385 762 387
rect 764 385 765 387
rect 841 499 842 501
rect 844 499 845 501
rect 841 505 842 507
rect 844 505 845 507
rect 941 559 942 561
rect 944 559 945 561
rect 941 565 942 567
rect 944 565 945 567
rect 1061 659 1062 661
rect 1064 659 1065 661
rect 1061 665 1062 667
rect 1064 665 1065 667
rect 601 719 602 721
rect 604 719 605 721
rect 601 725 602 727
rect 604 725 605 727
rect 441 519 442 521
rect 444 519 445 521
rect 441 525 442 527
rect 444 525 445 527
rect 741 759 742 761
rect 744 759 745 761
rect 741 765 742 767
rect 744 765 745 767
rect 341 559 342 561
rect 344 559 345 561
rect 341 565 342 567
rect 344 565 345 567
rect 361 559 362 561
rect 364 559 365 561
rect 361 565 362 567
rect 364 565 365 567
rect 821 399 822 401
rect 824 399 825 401
rect 821 405 822 407
rect 824 405 825 407
rect 641 1079 642 1081
rect 644 1079 645 1081
rect 641 1085 642 1087
rect 644 1085 645 1087
rect 681 519 682 521
rect 684 519 685 521
rect 681 525 682 527
rect 684 525 685 527
rect 761 639 762 641
rect 764 639 765 641
rect 761 645 762 647
rect 764 645 765 647
rect 821 819 822 821
rect 824 819 825 821
rect 821 825 822 827
rect 824 825 825 827
rect 761 419 762 421
rect 764 419 765 421
rect 761 425 762 427
rect 764 425 765 427
rect 501 879 502 881
rect 504 879 505 881
rect 501 885 502 887
rect 504 885 505 887
rect 621 599 622 601
rect 624 599 625 601
rect 621 605 622 607
rect 624 605 625 607
rect 261 699 262 701
rect 264 699 265 701
rect 261 705 262 707
rect 264 705 265 707
rect 801 499 802 501
rect 804 499 805 501
rect 801 505 802 507
rect 804 505 805 507
rect 421 799 422 801
rect 424 799 425 801
rect 421 805 422 807
rect 424 805 425 807
rect 861 439 862 441
rect 864 439 865 441
rect 861 445 862 447
rect 864 445 865 447
rect 761 1039 762 1041
rect 764 1039 765 1041
rect 761 1045 762 1047
rect 764 1045 765 1047
rect 821 919 822 921
rect 824 919 825 921
rect 821 925 822 927
rect 824 925 825 927
rect 681 779 682 781
rect 684 779 685 781
rect 681 785 682 787
rect 684 785 685 787
rect 661 499 662 501
rect 664 499 665 501
rect 661 505 662 507
rect 664 505 665 507
rect 721 979 722 981
rect 724 979 725 981
rect 721 985 722 987
rect 724 985 725 987
rect 581 659 582 661
rect 584 659 585 661
rect 581 665 582 667
rect 584 665 585 667
rect 941 759 942 761
rect 944 759 945 761
rect 941 765 942 767
rect 944 765 945 767
rect 861 539 862 541
rect 864 539 865 541
rect 861 545 862 547
rect 864 545 865 547
rect 1041 639 1042 641
rect 1044 639 1045 641
rect 1041 645 1042 647
rect 1044 645 1045 647
rect 701 819 702 821
rect 704 819 705 821
rect 701 825 702 827
rect 704 825 705 827
rect 821 859 822 861
rect 824 859 825 861
rect 821 865 822 867
rect 824 865 825 867
rect 961 619 962 621
rect 964 619 965 621
rect 961 625 962 627
rect 964 625 965 627
rect 541 379 542 381
rect 544 379 545 381
rect 541 385 542 387
rect 544 385 545 387
rect 701 939 702 941
rect 704 939 705 941
rect 701 945 702 947
rect 704 945 705 947
rect 641 659 642 661
rect 644 659 645 661
rect 641 665 642 667
rect 644 665 645 667
rect 701 879 702 881
rect 704 879 705 881
rect 701 885 702 887
rect 704 885 705 887
rect 661 539 662 541
rect 664 539 665 541
rect 661 545 662 547
rect 664 545 665 547
rect 741 679 742 681
rect 744 679 745 681
rect 741 685 742 687
rect 744 685 745 687
rect 621 339 622 341
rect 624 339 625 341
rect 621 345 622 347
rect 624 345 625 347
rect 881 579 882 581
rect 884 579 885 581
rect 881 585 882 587
rect 884 585 885 587
rect 701 759 702 761
rect 704 759 705 761
rect 701 765 702 767
rect 704 765 705 767
rect 701 719 702 721
rect 704 719 705 721
rect 701 725 702 727
rect 704 725 705 727
rect 601 559 602 561
rect 604 559 605 561
rect 601 565 602 567
rect 604 565 605 567
rect 581 1039 582 1041
rect 584 1039 585 1041
rect 581 1045 582 1047
rect 584 1045 585 1047
rect 721 539 722 541
rect 724 539 725 541
rect 721 545 722 547
rect 724 545 725 547
rect 621 519 622 521
rect 624 519 625 521
rect 621 525 622 527
rect 624 525 625 527
rect 641 779 642 781
rect 644 779 645 781
rect 641 785 642 787
rect 644 785 645 787
rect 521 579 522 581
rect 524 579 525 581
rect 521 585 522 587
rect 524 585 525 587
rect 521 659 522 661
rect 524 659 525 661
rect 521 665 522 667
rect 524 665 525 667
rect 801 859 802 861
rect 804 859 805 861
rect 801 865 802 867
rect 804 865 805 867
rect 321 599 322 601
rect 324 599 325 601
rect 321 605 322 607
rect 324 605 325 607
rect 541 459 542 461
rect 544 459 545 461
rect 541 465 542 467
rect 544 465 545 467
rect 801 899 802 901
rect 804 899 805 901
rect 801 905 802 907
rect 804 905 805 907
rect 601 999 602 1001
rect 604 999 605 1001
rect 601 1005 602 1007
rect 604 1005 605 1007
rect 441 859 442 861
rect 444 859 445 861
rect 441 865 442 867
rect 444 865 445 867
rect 721 419 722 421
rect 724 419 725 421
rect 721 425 722 427
rect 724 425 725 427
rect 581 719 582 721
rect 584 719 585 721
rect 581 725 582 727
rect 584 725 585 727
rect 741 659 742 661
rect 744 659 745 661
rect 741 665 742 667
rect 744 665 745 667
rect 821 619 822 621
rect 824 619 825 621
rect 821 625 822 627
rect 824 625 825 627
rect 361 719 362 721
rect 364 719 365 721
rect 361 725 362 727
rect 364 725 365 727
rect 541 939 542 941
rect 544 939 545 941
rect 541 945 542 947
rect 544 945 545 947
rect 541 679 542 681
rect 544 679 545 681
rect 541 685 542 687
rect 544 685 545 687
rect 961 639 962 641
rect 964 639 965 641
rect 961 645 962 647
rect 964 645 965 647
rect 581 839 582 841
rect 584 839 585 841
rect 581 845 582 847
rect 584 845 585 847
rect 721 899 722 901
rect 724 899 725 901
rect 721 905 722 907
rect 724 905 725 907
rect 661 839 662 841
rect 664 839 665 841
rect 661 845 662 847
rect 664 845 665 847
rect 701 299 702 301
rect 704 299 705 301
rect 701 305 702 307
rect 704 305 705 307
rect 441 759 442 761
rect 444 759 445 761
rect 441 765 442 767
rect 444 765 445 767
rect 441 539 442 541
rect 444 539 445 541
rect 441 545 442 547
rect 444 545 445 547
rect 461 459 462 461
rect 464 459 465 461
rect 461 465 462 467
rect 464 465 465 467
rect 401 699 402 701
rect 404 699 405 701
rect 401 705 402 707
rect 404 705 405 707
rect 681 479 682 481
rect 684 479 685 481
rect 681 485 682 487
rect 684 485 685 487
rect 681 339 682 341
rect 684 339 685 341
rect 681 345 682 347
rect 684 345 685 347
rect 721 919 722 921
rect 724 919 725 921
rect 721 925 722 927
rect 724 925 725 927
rect 541 859 542 861
rect 544 859 545 861
rect 541 865 542 867
rect 544 865 545 867
rect 701 1039 702 1041
rect 704 1039 705 1041
rect 701 1045 702 1047
rect 704 1045 705 1047
rect 781 979 782 981
rect 784 979 785 981
rect 781 985 782 987
rect 784 985 785 987
rect 921 519 922 521
rect 924 519 925 521
rect 921 525 922 527
rect 924 525 925 527
rect 461 599 462 601
rect 464 599 465 601
rect 461 605 462 607
rect 464 605 465 607
rect 861 679 862 681
rect 864 679 865 681
rect 861 685 862 687
rect 864 685 865 687
rect 661 739 662 741
rect 664 739 665 741
rect 661 745 662 747
rect 664 745 665 747
rect 481 579 482 581
rect 484 579 485 581
rect 481 585 482 587
rect 484 585 485 587
rect 821 639 822 641
rect 824 639 825 641
rect 821 645 822 647
rect 824 645 825 647
rect 321 739 322 741
rect 324 739 325 741
rect 321 745 322 747
rect 324 745 325 747
rect 641 899 642 901
rect 644 899 645 901
rect 641 905 642 907
rect 644 905 645 907
rect 661 959 662 961
rect 664 959 665 961
rect 661 965 662 967
rect 664 965 665 967
rect 601 539 602 541
rect 604 539 605 541
rect 601 545 602 547
rect 604 545 605 547
rect 441 459 442 461
rect 444 459 445 461
rect 441 465 442 467
rect 444 465 445 467
rect 681 359 682 361
rect 684 359 685 361
rect 681 365 682 367
rect 684 365 685 367
rect 821 659 822 661
rect 824 659 825 661
rect 821 665 822 667
rect 824 665 825 667
rect 741 859 742 861
rect 744 859 745 861
rect 741 865 742 867
rect 744 865 745 867
rect 621 299 622 301
rect 624 299 625 301
rect 621 305 622 307
rect 624 305 625 307
rect 741 579 742 581
rect 744 579 745 581
rect 741 585 742 587
rect 744 585 745 587
rect 841 659 842 661
rect 844 659 845 661
rect 841 665 842 667
rect 844 665 845 667
rect 241 639 242 641
rect 244 639 245 641
rect 241 645 242 647
rect 244 645 245 647
rect 801 599 802 601
rect 804 599 805 601
rect 801 605 802 607
rect 804 605 805 607
rect 741 739 742 741
rect 744 739 745 741
rect 741 745 742 747
rect 744 745 745 747
rect 681 539 682 541
rect 684 539 685 541
rect 681 545 682 547
rect 684 545 685 547
rect 981 719 982 721
rect 984 719 985 721
rect 981 725 982 727
rect 984 725 985 727
rect 1021 739 1022 741
rect 1024 739 1025 741
rect 1021 745 1022 747
rect 1024 745 1025 747
rect 461 419 462 421
rect 464 419 465 421
rect 461 425 462 427
rect 464 425 465 427
rect 501 399 502 401
rect 504 399 505 401
rect 501 405 502 407
rect 504 405 505 407
rect 401 719 402 721
rect 404 719 405 721
rect 401 725 402 727
rect 404 725 405 727
rect 941 839 942 841
rect 944 839 945 841
rect 941 845 942 847
rect 944 845 945 847
rect 721 379 722 381
rect 724 379 725 381
rect 721 385 722 387
rect 724 385 725 387
rect 301 619 302 621
rect 304 619 305 621
rect 301 625 302 627
rect 304 625 305 627
rect 701 419 702 421
rect 704 419 705 421
rect 701 425 702 427
rect 704 425 705 427
rect 521 799 522 801
rect 524 799 525 801
rect 521 805 522 807
rect 524 805 525 807
rect 521 479 522 481
rect 524 479 525 481
rect 521 485 522 487
rect 524 485 525 487
rect 1001 639 1002 641
rect 1004 639 1005 641
rect 1001 645 1002 647
rect 1004 645 1005 647
rect 461 579 462 581
rect 464 579 465 581
rect 461 585 462 587
rect 464 585 465 587
rect 621 699 622 701
rect 624 699 625 701
rect 621 705 622 707
rect 624 705 625 707
rect 921 739 922 741
rect 924 739 925 741
rect 921 745 922 747
rect 924 745 925 747
rect 561 439 562 441
rect 564 439 565 441
rect 561 445 562 447
rect 564 445 565 447
rect 641 1039 642 1041
rect 644 1039 645 1041
rect 641 1045 642 1047
rect 644 1045 645 1047
rect 841 419 842 421
rect 844 419 845 421
rect 841 425 842 427
rect 844 425 845 427
rect 421 819 422 821
rect 424 819 425 821
rect 421 825 422 827
rect 424 825 425 827
rect 841 699 842 701
rect 844 699 845 701
rect 841 705 842 707
rect 844 705 845 707
rect 601 779 602 781
rect 604 779 605 781
rect 601 785 602 787
rect 604 785 605 787
rect 1061 699 1062 701
rect 1064 699 1065 701
rect 1061 705 1062 707
rect 1064 705 1065 707
rect 721 1019 722 1021
rect 724 1019 725 1021
rect 721 1025 722 1027
rect 724 1025 725 1027
rect 661 1019 662 1021
rect 664 1019 665 1021
rect 661 1025 662 1027
rect 664 1025 665 1027
rect 421 759 422 761
rect 424 759 425 761
rect 421 765 422 767
rect 424 765 425 767
rect 401 799 402 801
rect 404 799 405 801
rect 401 805 402 807
rect 404 805 405 807
rect 501 479 502 481
rect 504 479 505 481
rect 501 485 502 487
rect 504 485 505 487
rect 581 739 582 741
rect 584 739 585 741
rect 581 745 582 747
rect 584 745 585 747
rect 721 999 722 1001
rect 724 999 725 1001
rect 721 1005 722 1007
rect 724 1005 725 1007
rect 661 519 662 521
rect 664 519 665 521
rect 661 525 662 527
rect 664 525 665 527
rect 801 619 802 621
rect 804 619 805 621
rect 801 625 802 627
rect 804 625 805 627
rect 721 759 722 761
rect 724 759 725 761
rect 721 765 722 767
rect 724 765 725 767
rect 701 499 702 501
rect 704 499 705 501
rect 701 505 702 507
rect 704 505 705 507
rect 521 979 522 981
rect 524 979 525 981
rect 521 985 522 987
rect 524 985 525 987
rect 621 659 622 661
rect 624 659 625 661
rect 621 665 622 667
rect 624 665 625 667
rect 341 539 342 541
rect 344 539 345 541
rect 341 545 342 547
rect 344 545 345 547
rect 601 499 602 501
rect 604 499 605 501
rect 601 505 602 507
rect 604 505 605 507
rect 941 719 942 721
rect 944 719 945 721
rect 941 725 942 727
rect 944 725 945 727
rect 701 839 702 841
rect 704 839 705 841
rect 701 845 702 847
rect 704 845 705 847
rect 921 659 922 661
rect 924 659 925 661
rect 921 665 922 667
rect 924 665 925 667
rect 841 519 842 521
rect 844 519 845 521
rect 841 525 842 527
rect 844 525 845 527
rect 821 759 822 761
rect 824 759 825 761
rect 821 765 822 767
rect 824 765 825 767
rect 881 819 882 821
rect 884 819 885 821
rect 881 825 882 827
rect 884 825 885 827
rect 461 779 462 781
rect 464 779 465 781
rect 461 785 462 787
rect 464 785 465 787
rect 441 439 442 441
rect 444 439 445 441
rect 441 445 442 447
rect 444 445 445 447
rect 521 619 522 621
rect 524 619 525 621
rect 521 625 522 627
rect 524 625 525 627
rect 441 499 442 501
rect 444 499 445 501
rect 441 505 442 507
rect 444 505 445 507
rect 901 799 902 801
rect 904 799 905 801
rect 901 805 902 807
rect 904 805 905 807
rect 761 459 762 461
rect 764 459 765 461
rect 761 465 762 467
rect 764 465 765 467
rect 961 819 962 821
rect 964 819 965 821
rect 961 825 962 827
rect 964 825 965 827
rect 461 759 462 761
rect 464 759 465 761
rect 461 765 462 767
rect 464 765 465 767
rect 921 619 922 621
rect 924 619 925 621
rect 921 625 922 627
rect 924 625 925 627
rect 481 919 482 921
rect 484 919 485 921
rect 481 925 482 927
rect 484 925 485 927
rect 641 939 642 941
rect 644 939 645 941
rect 641 945 642 947
rect 644 945 645 947
rect 881 699 882 701
rect 884 699 885 701
rect 881 705 882 707
rect 884 705 885 707
rect 601 759 602 761
rect 604 759 605 761
rect 601 765 602 767
rect 604 765 605 767
rect 361 699 362 701
rect 364 699 365 701
rect 361 705 362 707
rect 364 705 365 707
rect 781 499 782 501
rect 784 499 785 501
rect 781 505 782 507
rect 784 505 785 507
rect 281 659 282 661
rect 284 659 285 661
rect 281 665 282 667
rect 284 665 285 667
rect 361 739 362 741
rect 364 739 365 741
rect 361 745 362 747
rect 364 745 365 747
rect 521 779 522 781
rect 524 779 525 781
rect 521 785 522 787
rect 524 785 525 787
rect 401 479 402 481
rect 404 479 405 481
rect 401 485 402 487
rect 404 485 405 487
rect 541 779 542 781
rect 544 779 545 781
rect 541 785 542 787
rect 544 785 545 787
rect 401 739 402 741
rect 404 739 405 741
rect 401 745 402 747
rect 404 745 405 747
rect 561 939 562 941
rect 564 939 565 941
rect 561 945 562 947
rect 564 945 565 947
rect 861 819 862 821
rect 864 819 865 821
rect 861 825 862 827
rect 864 825 865 827
rect 681 619 682 621
rect 684 619 685 621
rect 681 625 682 627
rect 684 625 685 627
rect 901 719 902 721
rect 904 719 905 721
rect 901 725 902 727
rect 904 725 905 727
rect 781 919 782 921
rect 784 919 785 921
rect 781 925 782 927
rect 784 925 785 927
rect 741 939 742 941
rect 744 939 745 941
rect 741 945 742 947
rect 744 945 745 947
rect 1001 659 1002 661
rect 1004 659 1005 661
rect 1001 665 1002 667
rect 1004 665 1005 667
rect 761 339 762 341
rect 764 339 765 341
rect 761 345 762 347
rect 764 345 765 347
rect 681 319 682 321
rect 684 319 685 321
rect 681 325 682 327
rect 684 325 685 327
rect 621 539 622 541
rect 624 539 625 541
rect 621 545 622 547
rect 624 545 625 547
rect 501 559 502 561
rect 504 559 505 561
rect 501 565 502 567
rect 504 565 505 567
rect 961 739 962 741
rect 964 739 965 741
rect 961 745 962 747
rect 964 745 965 747
rect 381 839 382 841
rect 384 839 385 841
rect 381 845 382 847
rect 384 845 385 847
rect 661 579 662 581
rect 664 579 665 581
rect 661 585 662 587
rect 664 585 665 587
rect 621 739 622 741
rect 624 739 625 741
rect 621 745 622 747
rect 624 745 625 747
rect 701 659 702 661
rect 704 659 705 661
rect 701 665 702 667
rect 704 665 705 667
rect 321 659 322 661
rect 324 659 325 661
rect 321 665 322 667
rect 324 665 325 667
rect 321 719 322 721
rect 324 719 325 721
rect 321 725 322 727
rect 324 725 325 727
rect 1041 679 1042 681
rect 1044 679 1045 681
rect 1041 685 1042 687
rect 1044 685 1045 687
rect 541 899 542 901
rect 544 899 545 901
rect 541 905 542 907
rect 544 905 545 907
rect 881 519 882 521
rect 884 519 885 521
rect 881 525 882 527
rect 884 525 885 527
rect 301 639 302 641
rect 304 639 305 641
rect 301 645 302 647
rect 304 645 305 647
rect 421 779 422 781
rect 424 779 425 781
rect 421 785 422 787
rect 424 785 425 787
rect 641 859 642 861
rect 644 859 645 861
rect 641 865 642 867
rect 644 865 645 867
rect 881 499 882 501
rect 884 499 885 501
rect 881 505 882 507
rect 884 505 885 507
rect 401 819 402 821
rect 404 819 405 821
rect 401 825 402 827
rect 404 825 405 827
rect 841 819 842 821
rect 844 819 845 821
rect 841 825 842 827
rect 844 825 845 827
rect 541 399 542 401
rect 544 399 545 401
rect 541 405 542 407
rect 544 405 545 407
rect 541 419 542 421
rect 544 419 545 421
rect 541 425 542 427
rect 544 425 545 427
rect 841 539 842 541
rect 844 539 845 541
rect 841 545 842 547
rect 844 545 845 547
rect 981 799 982 801
rect 984 799 985 801
rect 981 805 982 807
rect 984 805 985 807
rect 521 399 522 401
rect 524 399 525 401
rect 521 405 522 407
rect 524 405 525 407
rect 861 659 862 661
rect 864 659 865 661
rect 861 665 862 667
rect 864 665 865 667
rect 581 319 582 321
rect 584 319 585 321
rect 581 325 582 327
rect 584 325 585 327
rect 761 559 762 561
rect 764 559 765 561
rect 761 565 762 567
rect 764 565 765 567
rect 901 779 902 781
rect 904 779 905 781
rect 901 785 902 787
rect 904 785 905 787
rect 981 619 982 621
rect 984 619 985 621
rect 981 625 982 627
rect 984 625 985 627
rect 681 559 682 561
rect 684 559 685 561
rect 681 565 682 567
rect 684 565 685 567
rect 881 459 882 461
rect 884 459 885 461
rect 881 465 882 467
rect 884 465 885 467
rect 761 839 762 841
rect 764 839 765 841
rect 761 845 762 847
rect 764 845 765 847
rect 921 599 922 601
rect 924 599 925 601
rect 921 605 922 607
rect 924 605 925 607
rect 881 619 882 621
rect 884 619 885 621
rect 881 625 882 627
rect 884 625 885 627
rect 301 739 302 741
rect 304 739 305 741
rect 301 745 302 747
rect 304 745 305 747
rect 1021 659 1022 661
rect 1024 659 1025 661
rect 1021 665 1022 667
rect 1024 665 1025 667
rect 661 979 662 981
rect 664 979 665 981
rect 661 985 662 987
rect 664 985 665 987
rect 801 419 802 421
rect 804 419 805 421
rect 801 425 802 427
rect 804 425 805 427
rect 1001 599 1002 601
rect 1004 599 1005 601
rect 1001 605 1002 607
rect 1004 605 1005 607
rect 861 559 862 561
rect 864 559 865 561
rect 861 565 862 567
rect 864 565 865 567
rect 381 699 382 701
rect 384 699 385 701
rect 381 705 382 707
rect 384 705 385 707
rect 661 659 662 661
rect 664 659 665 661
rect 661 665 662 667
rect 664 665 665 667
rect 521 939 522 941
rect 524 939 525 941
rect 521 945 522 947
rect 524 945 525 947
rect 741 799 742 801
rect 744 799 745 801
rect 741 805 742 807
rect 744 805 745 807
rect 521 499 522 501
rect 524 499 525 501
rect 521 505 522 507
rect 524 505 525 507
rect 541 479 542 481
rect 544 479 545 481
rect 541 485 542 487
rect 544 485 545 487
rect 401 579 402 581
rect 404 579 405 581
rect 401 585 402 587
rect 404 585 405 587
rect 981 639 982 641
rect 984 639 985 641
rect 981 645 982 647
rect 984 645 985 647
rect 461 819 462 821
rect 464 819 465 821
rect 461 825 462 827
rect 464 825 465 827
rect 581 479 582 481
rect 584 479 585 481
rect 581 485 582 487
rect 584 485 585 487
rect 421 579 422 581
rect 424 579 425 581
rect 421 585 422 587
rect 424 585 425 587
rect 401 779 402 781
rect 404 779 405 781
rect 401 785 402 787
rect 404 785 405 787
rect 301 799 302 801
rect 304 799 305 801
rect 301 805 302 807
rect 304 805 305 807
rect 941 519 942 521
rect 944 519 945 521
rect 941 525 942 527
rect 944 525 945 527
rect 581 999 582 1001
rect 584 999 585 1001
rect 581 1005 582 1007
rect 584 1005 585 1007
rect 681 279 682 281
rect 684 279 685 281
rect 681 285 682 287
rect 684 285 685 287
rect 881 439 882 441
rect 884 439 885 441
rect 881 445 882 447
rect 884 445 885 447
rect 401 599 402 601
rect 404 599 405 601
rect 401 605 402 607
rect 404 605 405 607
rect 901 559 902 561
rect 904 559 905 561
rect 901 565 902 567
rect 904 565 905 567
rect 1001 759 1002 761
rect 1004 759 1005 761
rect 1001 765 1002 767
rect 1004 765 1005 767
rect 321 639 322 641
rect 324 639 325 641
rect 321 645 322 647
rect 324 645 325 647
rect 681 879 682 881
rect 684 879 685 881
rect 681 885 682 887
rect 684 885 685 887
rect 861 799 862 801
rect 864 799 865 801
rect 861 805 862 807
rect 864 805 865 807
rect 861 699 862 701
rect 864 699 865 701
rect 861 705 862 707
rect 864 705 865 707
rect 1001 679 1002 681
rect 1004 679 1005 681
rect 1001 685 1002 687
rect 1004 685 1005 687
rect 741 699 742 701
rect 744 699 745 701
rect 741 705 742 707
rect 744 705 745 707
rect 301 679 302 681
rect 304 679 305 681
rect 301 685 302 687
rect 304 685 305 687
rect 681 759 682 761
rect 684 759 685 761
rect 681 765 682 767
rect 684 765 685 767
rect 661 399 662 401
rect 664 399 665 401
rect 661 405 662 407
rect 664 405 665 407
rect 381 719 382 721
rect 384 719 385 721
rect 381 725 382 727
rect 384 725 385 727
rect 301 719 302 721
rect 304 719 305 721
rect 301 725 302 727
rect 304 725 305 727
rect 701 979 702 981
rect 704 979 705 981
rect 701 985 702 987
rect 704 985 705 987
rect 541 739 542 741
rect 544 739 545 741
rect 541 745 542 747
rect 544 745 545 747
rect 821 719 822 721
rect 824 719 825 721
rect 821 725 822 727
rect 824 725 825 727
rect 641 759 642 761
rect 644 759 645 761
rect 641 765 642 767
rect 644 765 645 767
rect 761 599 762 601
rect 764 599 765 601
rect 761 605 762 607
rect 764 605 765 607
rect 841 579 842 581
rect 844 579 845 581
rect 841 585 842 587
rect 844 585 845 587
rect 421 599 422 601
rect 424 599 425 601
rect 421 605 422 607
rect 424 605 425 607
rect 741 439 742 441
rect 744 439 745 441
rect 741 445 742 447
rect 744 445 745 447
rect 801 959 802 961
rect 804 959 805 961
rect 801 965 802 967
rect 804 965 805 967
rect 781 859 782 861
rect 784 859 785 861
rect 781 865 782 867
rect 784 865 785 867
rect 681 1019 682 1021
rect 684 1019 685 1021
rect 681 1025 682 1027
rect 684 1025 685 1027
rect 541 959 542 961
rect 544 959 545 961
rect 541 965 542 967
rect 544 965 545 967
rect 981 599 982 601
rect 984 599 985 601
rect 981 605 982 607
rect 984 605 985 607
rect 801 919 802 921
rect 804 919 805 921
rect 801 925 802 927
rect 804 925 805 927
rect 961 659 962 661
rect 964 659 965 661
rect 961 665 962 667
rect 964 665 965 667
rect 641 999 642 1001
rect 644 999 645 1001
rect 641 1005 642 1007
rect 644 1005 645 1007
rect 321 579 322 581
rect 324 579 325 581
rect 321 585 322 587
rect 324 585 325 587
rect 581 339 582 341
rect 584 339 585 341
rect 581 345 582 347
rect 584 345 585 347
rect 581 819 582 821
rect 584 819 585 821
rect 581 825 582 827
rect 584 825 585 827
rect 761 819 762 821
rect 764 819 765 821
rect 761 825 762 827
rect 764 825 765 827
rect 581 859 582 861
rect 584 859 585 861
rect 581 865 582 867
rect 584 865 585 867
rect 701 619 702 621
rect 704 619 705 621
rect 701 625 702 627
rect 704 625 705 627
rect 521 599 522 601
rect 524 599 525 601
rect 521 605 522 607
rect 524 605 525 607
rect 581 919 582 921
rect 584 919 585 921
rect 581 925 582 927
rect 584 925 585 927
rect 881 659 882 661
rect 884 659 885 661
rect 881 665 882 667
rect 884 665 885 667
rect 461 879 462 881
rect 464 879 465 881
rect 461 885 462 887
rect 464 885 465 887
rect 521 899 522 901
rect 524 899 525 901
rect 521 905 522 907
rect 524 905 525 907
rect 881 679 882 681
rect 884 679 885 681
rect 881 685 882 687
rect 884 685 885 687
rect 441 779 442 781
rect 444 779 445 781
rect 441 785 442 787
rect 444 785 445 787
rect 401 859 402 861
rect 404 859 405 861
rect 401 865 402 867
rect 404 865 405 867
rect 681 959 682 961
rect 684 959 685 961
rect 681 965 682 967
rect 684 965 685 967
rect 821 459 822 461
rect 824 459 825 461
rect 821 465 822 467
rect 824 465 825 467
rect 721 499 722 501
rect 724 499 725 501
rect 721 505 722 507
rect 724 505 725 507
rect 501 819 502 821
rect 504 819 505 821
rect 501 825 502 827
rect 504 825 505 827
rect 441 799 442 801
rect 444 799 445 801
rect 441 805 442 807
rect 444 805 445 807
rect 761 739 762 741
rect 764 739 765 741
rect 761 745 762 747
rect 764 745 765 747
rect 901 659 902 661
rect 904 659 905 661
rect 901 665 902 667
rect 904 665 905 667
rect 561 799 562 801
rect 564 799 565 801
rect 561 805 562 807
rect 564 805 565 807
rect 921 819 922 821
rect 924 819 925 821
rect 921 825 922 827
rect 924 825 925 827
rect 381 739 382 741
rect 384 739 385 741
rect 381 745 382 747
rect 384 745 385 747
rect 661 699 662 701
rect 664 699 665 701
rect 661 705 662 707
rect 664 705 665 707
rect 541 839 542 841
rect 544 839 545 841
rect 541 845 542 847
rect 544 845 545 847
rect 301 579 302 581
rect 304 579 305 581
rect 301 585 302 587
rect 304 585 305 587
rect 781 699 782 701
rect 784 699 785 701
rect 781 705 782 707
rect 784 705 785 707
rect 481 899 482 901
rect 484 899 485 901
rect 481 905 482 907
rect 484 905 485 907
rect 741 999 742 1001
rect 744 999 745 1001
rect 741 1005 742 1007
rect 744 1005 745 1007
rect 661 479 662 481
rect 664 479 665 481
rect 661 485 662 487
rect 664 485 665 487
rect 481 719 482 721
rect 484 719 485 721
rect 481 725 482 727
rect 484 725 485 727
rect 861 579 862 581
rect 864 579 865 581
rect 861 585 862 587
rect 864 585 865 587
rect 421 499 422 501
rect 424 499 425 501
rect 421 505 422 507
rect 424 505 425 507
rect 501 499 502 501
rect 504 499 505 501
rect 501 505 502 507
rect 504 505 505 507
rect 641 679 642 681
rect 644 679 645 681
rect 641 685 642 687
rect 644 685 645 687
rect 901 739 902 741
rect 904 739 905 741
rect 901 745 902 747
rect 904 745 905 747
rect 601 959 602 961
rect 604 959 605 961
rect 601 965 602 967
rect 604 965 605 967
rect 661 719 662 721
rect 664 719 665 721
rect 661 725 662 727
rect 664 725 665 727
rect 781 799 782 801
rect 784 799 785 801
rect 781 805 782 807
rect 784 805 785 807
rect 841 759 842 761
rect 844 759 845 761
rect 841 765 842 767
rect 844 765 845 767
rect 621 819 622 821
rect 624 819 625 821
rect 621 825 622 827
rect 624 825 625 827
rect 381 659 382 661
rect 384 659 385 661
rect 381 665 382 667
rect 384 665 385 667
rect 721 699 722 701
rect 724 699 725 701
rect 721 705 722 707
rect 724 705 725 707
rect 761 759 762 761
rect 764 759 765 761
rect 761 765 762 767
rect 764 765 765 767
rect 641 439 642 441
rect 644 439 645 441
rect 641 445 642 447
rect 644 445 645 447
rect 821 419 822 421
rect 824 419 825 421
rect 821 425 822 427
rect 824 425 825 427
rect 441 659 442 661
rect 444 659 445 661
rect 441 665 442 667
rect 444 665 445 667
rect 781 619 782 621
rect 784 619 785 621
rect 781 625 782 627
rect 784 625 785 627
rect 281 679 282 681
rect 284 679 285 681
rect 281 685 282 687
rect 284 685 285 687
rect 741 919 742 921
rect 744 919 745 921
rect 741 925 742 927
rect 744 925 745 927
rect 421 559 422 561
rect 424 559 425 561
rect 421 565 422 567
rect 424 565 425 567
rect 461 799 462 801
rect 464 799 465 801
rect 461 805 462 807
rect 464 805 465 807
rect 461 479 462 481
rect 464 479 465 481
rect 461 485 462 487
rect 464 485 465 487
rect 841 639 842 641
rect 844 639 845 641
rect 841 645 842 647
rect 844 645 845 647
rect 361 779 362 781
rect 364 779 365 781
rect 361 785 362 787
rect 364 785 365 787
rect 621 939 622 941
rect 624 939 625 941
rect 621 945 622 947
rect 624 945 625 947
rect 881 739 882 741
rect 884 739 885 741
rect 881 745 882 747
rect 884 745 885 747
rect 821 939 822 941
rect 824 939 825 941
rect 821 945 822 947
rect 824 945 825 947
rect 601 859 602 861
rect 604 859 605 861
rect 601 865 602 867
rect 604 865 605 867
rect 681 819 682 821
rect 684 819 685 821
rect 681 825 682 827
rect 684 825 685 827
rect 821 579 822 581
rect 824 579 825 581
rect 821 585 822 587
rect 824 585 825 587
rect 621 619 622 621
rect 624 619 625 621
rect 621 625 622 627
rect 624 625 625 627
rect 601 879 602 881
rect 604 879 605 881
rect 601 885 602 887
rect 604 885 605 887
rect 381 499 382 501
rect 384 499 385 501
rect 381 505 382 507
rect 384 505 385 507
rect 581 499 582 501
rect 584 499 585 501
rect 581 505 582 507
rect 584 505 585 507
rect 881 799 882 801
rect 884 799 885 801
rect 881 805 882 807
rect 884 805 885 807
rect 581 519 582 521
rect 584 519 585 521
rect 581 525 582 527
rect 584 525 585 527
rect 881 779 882 781
rect 884 779 885 781
rect 881 785 882 787
rect 884 785 885 787
rect 521 379 522 381
rect 524 379 525 381
rect 521 385 522 387
rect 524 385 525 387
rect 881 879 882 881
rect 884 879 885 881
rect 881 885 882 887
rect 884 885 885 887
rect 461 699 462 701
rect 464 699 465 701
rect 461 705 462 707
rect 464 705 465 707
rect 281 639 282 641
rect 284 639 285 641
rect 281 645 282 647
rect 284 645 285 647
rect 701 439 702 441
rect 704 439 705 441
rect 701 445 702 447
rect 704 445 705 447
rect 641 359 642 361
rect 644 359 645 361
rect 641 365 642 367
rect 644 365 645 367
rect 861 719 862 721
rect 864 719 865 721
rect 861 725 862 727
rect 864 725 865 727
rect 961 779 962 781
rect 964 779 965 781
rect 961 785 962 787
rect 964 785 965 787
rect 1021 719 1022 721
rect 1024 719 1025 721
rect 1021 725 1022 727
rect 1024 725 1025 727
rect 881 839 882 841
rect 884 839 885 841
rect 881 845 882 847
rect 884 845 885 847
rect 641 419 642 421
rect 644 419 645 421
rect 641 425 642 427
rect 644 425 645 427
rect 841 599 842 601
rect 844 599 845 601
rect 841 605 842 607
rect 844 605 845 607
rect 561 559 562 561
rect 564 559 565 561
rect 561 565 562 567
rect 564 565 565 567
rect 741 899 742 901
rect 744 899 745 901
rect 741 905 742 907
rect 744 905 745 907
rect 581 959 582 961
rect 584 959 585 961
rect 581 965 582 967
rect 584 965 585 967
rect 501 899 502 901
rect 504 899 505 901
rect 501 905 502 907
rect 504 905 505 907
rect 461 519 462 521
rect 464 519 465 521
rect 461 525 462 527
rect 464 525 465 527
rect 681 579 682 581
rect 684 579 685 581
rect 681 585 682 587
rect 684 585 685 587
rect 941 679 942 681
rect 944 679 945 681
rect 941 685 942 687
rect 944 685 945 687
rect 901 519 902 521
rect 904 519 905 521
rect 901 525 902 527
rect 904 525 905 527
rect 601 399 602 401
rect 604 399 605 401
rect 601 405 602 407
rect 604 405 605 407
rect 581 439 582 441
rect 584 439 585 441
rect 581 445 582 447
rect 584 445 585 447
rect 561 499 562 501
rect 564 499 565 501
rect 561 505 562 507
rect 564 505 565 507
rect 501 859 502 861
rect 504 859 505 861
rect 501 865 502 867
rect 504 865 505 867
rect 481 819 482 821
rect 484 819 485 821
rect 481 825 482 827
rect 484 825 485 827
rect 721 859 722 861
rect 724 859 725 861
rect 721 865 722 867
rect 724 865 725 867
rect 601 439 602 441
rect 604 439 605 441
rect 601 445 602 447
rect 604 445 605 447
rect 821 539 822 541
rect 824 539 825 541
rect 821 545 822 547
rect 824 545 825 547
rect 661 359 662 361
rect 664 359 665 361
rect 661 365 662 367
rect 664 365 665 367
rect 581 759 582 761
rect 584 759 585 761
rect 581 765 582 767
rect 584 765 585 767
rect 601 939 602 941
rect 604 939 605 941
rect 601 945 602 947
rect 604 945 605 947
rect 521 699 522 701
rect 524 699 525 701
rect 521 705 522 707
rect 524 705 525 707
rect 681 499 682 501
rect 684 499 685 501
rect 681 505 682 507
rect 684 505 685 507
rect 781 679 782 681
rect 784 679 785 681
rect 781 685 782 687
rect 784 685 785 687
rect 281 599 282 601
rect 284 599 285 601
rect 281 605 282 607
rect 284 605 285 607
rect 681 939 682 941
rect 684 939 685 941
rect 681 945 682 947
rect 684 945 685 947
rect 261 619 262 621
rect 264 619 265 621
rect 261 625 262 627
rect 264 625 265 627
rect 701 539 702 541
rect 704 539 705 541
rect 701 545 702 547
rect 704 545 705 547
rect 641 499 642 501
rect 644 499 645 501
rect 641 505 642 507
rect 644 505 645 507
rect 901 699 902 701
rect 904 699 905 701
rect 901 705 902 707
rect 904 705 905 707
rect 501 679 502 681
rect 504 679 505 681
rect 501 685 502 687
rect 504 685 505 687
rect 481 939 482 941
rect 484 939 485 941
rect 481 945 482 947
rect 484 945 485 947
rect 661 339 662 341
rect 664 339 665 341
rect 661 345 662 347
rect 664 345 665 347
rect 441 739 442 741
rect 444 739 445 741
rect 441 745 442 747
rect 444 745 445 747
rect 721 839 722 841
rect 724 839 725 841
rect 721 845 722 847
rect 724 845 725 847
rect 701 859 702 861
rect 704 859 705 861
rect 701 865 702 867
rect 704 865 705 867
rect 461 439 462 441
rect 464 439 465 441
rect 461 445 462 447
rect 464 445 465 447
rect 741 339 742 341
rect 744 339 745 341
rect 741 345 742 347
rect 744 345 745 347
rect 461 1039 462 1041
rect 464 1039 465 1041
rect 461 1045 462 1047
rect 464 1045 465 1047
rect 641 299 642 301
rect 644 299 645 301
rect 641 305 642 307
rect 644 305 645 307
rect 1041 659 1042 661
rect 1044 659 1045 661
rect 1041 665 1042 667
rect 1044 665 1045 667
rect 501 419 502 421
rect 504 419 505 421
rect 501 425 502 427
rect 504 425 505 427
rect 681 799 682 801
rect 684 799 685 801
rect 681 805 682 807
rect 684 805 685 807
rect 721 619 722 621
rect 724 619 725 621
rect 721 625 722 627
rect 724 625 725 627
rect 341 619 342 621
rect 344 619 345 621
rect 341 625 342 627
rect 344 625 345 627
rect 421 639 422 641
rect 424 639 425 641
rect 421 645 422 647
rect 424 645 425 647
rect 821 379 822 381
rect 824 379 825 381
rect 821 385 822 387
rect 824 385 825 387
rect 361 519 362 521
rect 364 519 365 521
rect 361 525 362 527
rect 364 525 365 527
rect 441 819 442 821
rect 444 819 445 821
rect 441 825 442 827
rect 444 825 445 827
rect 561 919 562 921
rect 564 919 565 921
rect 561 925 562 927
rect 564 925 565 927
rect 821 739 822 741
rect 824 739 825 741
rect 821 745 822 747
rect 824 745 825 747
rect 921 759 922 761
rect 924 759 925 761
rect 921 765 922 767
rect 924 765 925 767
rect 621 859 622 861
rect 624 859 625 861
rect 621 865 622 867
rect 624 865 625 867
rect 681 379 682 381
rect 684 379 685 381
rect 681 385 682 387
rect 684 385 685 387
rect 701 559 702 561
rect 704 559 705 561
rect 701 565 702 567
rect 704 565 705 567
rect 921 499 922 501
rect 924 499 925 501
rect 921 505 922 507
rect 924 505 925 507
rect 541 439 542 441
rect 544 439 545 441
rect 541 445 542 447
rect 544 445 545 447
rect 501 539 502 541
rect 504 539 505 541
rect 501 545 502 547
rect 504 545 505 547
rect 941 739 942 741
rect 944 739 945 741
rect 941 745 942 747
rect 944 745 945 747
rect 841 859 842 861
rect 844 859 845 861
rect 841 865 842 867
rect 844 865 845 867
rect 821 439 822 441
rect 824 439 825 441
rect 821 445 822 447
rect 824 445 825 447
rect 941 639 942 641
rect 944 639 945 641
rect 941 645 942 647
rect 944 645 945 647
rect 521 459 522 461
rect 524 459 525 461
rect 521 465 522 467
rect 524 465 525 467
rect 1001 739 1002 741
rect 1004 739 1005 741
rect 1001 745 1002 747
rect 1004 745 1005 747
rect 681 999 682 1001
rect 684 999 685 1001
rect 681 1005 682 1007
rect 684 1005 685 1007
rect 501 639 502 641
rect 504 639 505 641
rect 501 645 502 647
rect 504 645 505 647
rect 961 719 962 721
rect 964 719 965 721
rect 961 725 962 727
rect 964 725 965 727
rect 701 599 702 601
rect 704 599 705 601
rect 701 605 702 607
rect 704 605 705 607
rect 581 559 582 561
rect 584 559 585 561
rect 581 565 582 567
rect 584 565 585 567
rect 761 899 762 901
rect 764 899 765 901
rect 761 905 762 907
rect 764 905 765 907
rect 761 859 762 861
rect 764 859 765 861
rect 761 865 762 867
rect 764 865 765 867
rect 601 659 602 661
rect 604 659 605 661
rect 601 665 602 667
rect 604 665 605 667
rect 861 619 862 621
rect 864 619 865 621
rect 861 625 862 627
rect 864 625 865 627
rect 901 499 902 501
rect 904 499 905 501
rect 901 505 902 507
rect 904 505 905 507
rect 541 599 542 601
rect 544 599 545 601
rect 541 605 542 607
rect 544 605 545 607
rect 681 419 682 421
rect 684 419 685 421
rect 681 425 682 427
rect 684 425 685 427
rect 321 559 322 561
rect 324 559 325 561
rect 321 565 322 567
rect 324 565 325 567
rect 561 899 562 901
rect 564 899 565 901
rect 561 905 562 907
rect 564 905 565 907
rect 1021 679 1022 681
rect 1024 679 1025 681
rect 1021 685 1022 687
rect 1024 685 1025 687
rect 481 599 482 601
rect 484 599 485 601
rect 481 605 482 607
rect 484 605 485 607
rect 861 519 862 521
rect 864 519 865 521
rect 861 525 862 527
rect 864 525 865 527
rect 741 779 742 781
rect 744 779 745 781
rect 741 785 742 787
rect 744 785 745 787
rect 1041 699 1042 701
rect 1044 699 1045 701
rect 1041 705 1042 707
rect 1044 705 1045 707
rect 881 719 882 721
rect 884 719 885 721
rect 881 725 882 727
rect 884 725 885 727
rect 561 759 562 761
rect 564 759 565 761
rect 561 765 562 767
rect 564 765 565 767
rect 821 499 822 501
rect 824 499 825 501
rect 821 505 822 507
rect 824 505 825 507
rect 641 319 642 321
rect 644 319 645 321
rect 641 325 642 327
rect 644 325 645 327
rect 761 799 762 801
rect 764 799 765 801
rect 761 805 762 807
rect 764 805 765 807
rect 681 1039 682 1041
rect 684 1039 685 1041
rect 681 1045 682 1047
rect 684 1045 685 1047
rect 641 919 642 921
rect 644 919 645 921
rect 641 925 642 927
rect 644 925 645 927
rect 881 539 882 541
rect 884 539 885 541
rect 881 545 882 547
rect 884 545 885 547
rect 621 799 622 801
rect 624 799 625 801
rect 621 805 622 807
rect 624 805 625 807
rect 381 519 382 521
rect 384 519 385 521
rect 381 525 382 527
rect 384 525 385 527
rect 581 619 582 621
rect 584 619 585 621
rect 581 625 582 627
rect 584 625 585 627
rect 961 599 962 601
rect 964 599 965 601
rect 961 605 962 607
rect 964 605 965 607
rect 741 479 742 481
rect 744 479 745 481
rect 741 485 742 487
rect 744 485 745 487
rect 801 579 802 581
rect 804 579 805 581
rect 801 585 802 587
rect 804 585 805 587
rect 421 459 422 461
rect 424 459 425 461
rect 421 465 422 467
rect 424 465 425 467
rect 501 459 502 461
rect 504 459 505 461
rect 501 465 502 467
rect 504 465 505 467
rect 721 779 722 781
rect 724 779 725 781
rect 721 785 722 787
rect 724 785 725 787
rect 581 939 582 941
rect 584 939 585 941
rect 581 945 582 947
rect 584 945 585 947
rect 641 379 642 381
rect 644 379 645 381
rect 641 385 642 387
rect 644 385 645 387
rect 901 639 902 641
rect 904 639 905 641
rect 901 645 902 647
rect 904 645 905 647
rect 781 819 782 821
rect 784 819 785 821
rect 781 825 782 827
rect 784 825 785 827
rect 341 819 342 821
rect 344 819 345 821
rect 341 825 342 827
rect 344 825 345 827
rect 621 279 622 281
rect 624 279 625 281
rect 621 285 622 287
rect 624 285 625 287
rect 581 359 582 361
rect 584 359 585 361
rect 581 365 582 367
rect 584 365 585 367
rect 801 739 802 741
rect 804 739 805 741
rect 801 745 802 747
rect 804 745 805 747
rect 741 819 742 821
rect 744 819 745 821
rect 741 825 742 827
rect 744 825 745 827
rect 241 699 242 701
rect 244 699 245 701
rect 241 705 242 707
rect 244 705 245 707
rect 461 679 462 681
rect 464 679 465 681
rect 461 685 462 687
rect 464 685 465 687
rect 941 699 942 701
rect 944 699 945 701
rect 941 705 942 707
rect 944 705 945 707
rect 761 919 762 921
rect 764 919 765 921
rect 761 925 762 927
rect 764 925 765 927
rect 801 839 802 841
rect 804 839 805 841
rect 801 845 802 847
rect 804 845 805 847
rect 601 359 602 361
rect 604 359 605 361
rect 601 365 602 367
rect 604 365 605 367
rect 821 519 822 521
rect 824 519 825 521
rect 821 525 822 527
rect 824 525 825 527
rect 841 799 842 801
rect 844 799 845 801
rect 841 805 842 807
rect 844 805 845 807
rect 521 719 522 721
rect 524 719 525 721
rect 521 725 522 727
rect 524 725 525 727
rect 361 619 362 621
rect 364 619 365 621
rect 361 625 362 627
rect 364 625 365 627
rect 701 639 702 641
rect 704 639 705 641
rect 701 645 702 647
rect 704 645 705 647
rect 461 839 462 841
rect 464 839 465 841
rect 461 845 462 847
rect 464 845 465 847
rect 361 659 362 661
rect 364 659 365 661
rect 361 665 362 667
rect 364 665 365 667
rect 721 319 722 321
rect 724 319 725 321
rect 721 325 722 327
rect 724 325 725 327
rect 341 639 342 641
rect 344 639 345 641
rect 341 645 342 647
rect 344 645 345 647
rect 401 679 402 681
rect 404 679 405 681
rect 401 685 402 687
rect 404 685 405 687
rect 981 579 982 581
rect 984 579 985 581
rect 981 585 982 587
rect 984 585 985 587
rect 561 1019 562 1021
rect 564 1019 565 1021
rect 561 1025 562 1027
rect 564 1025 565 1027
rect 781 419 782 421
rect 784 419 785 421
rect 781 425 782 427
rect 784 425 785 427
rect 801 399 802 401
rect 804 399 805 401
rect 801 405 802 407
rect 804 405 805 407
rect 661 379 662 381
rect 664 379 665 381
rect 661 385 662 387
rect 664 385 665 387
rect 401 539 402 541
rect 404 539 405 541
rect 401 545 402 547
rect 404 545 405 547
rect 401 519 402 521
rect 404 519 405 521
rect 401 525 402 527
rect 404 525 405 527
rect 421 699 422 701
rect 424 699 425 701
rect 421 705 422 707
rect 424 705 425 707
rect 861 899 862 901
rect 864 899 865 901
rect 861 905 862 907
rect 864 905 865 907
rect 521 879 522 881
rect 524 879 525 881
rect 521 885 522 887
rect 524 885 525 887
rect 821 679 822 681
rect 824 679 825 681
rect 821 685 822 687
rect 824 685 825 687
rect 861 879 862 881
rect 864 879 865 881
rect 861 885 862 887
rect 864 885 865 887
rect 941 799 942 801
rect 944 799 945 801
rect 941 805 942 807
rect 944 805 945 807
rect 581 979 582 981
rect 584 979 585 981
rect 581 985 582 987
rect 584 985 585 987
rect 621 359 622 361
rect 624 359 625 361
rect 621 365 622 367
rect 624 365 625 367
rect 981 659 982 661
rect 984 659 985 661
rect 981 665 982 667
rect 984 665 985 667
rect 861 859 862 861
rect 864 859 865 861
rect 861 865 862 867
rect 864 865 865 867
rect 661 939 662 941
rect 664 939 665 941
rect 661 945 662 947
rect 664 945 665 947
rect 721 879 722 881
rect 724 879 725 881
rect 721 885 722 887
rect 724 885 725 887
rect 821 799 822 801
rect 824 799 825 801
rect 821 805 822 807
rect 824 805 825 807
rect 761 979 762 981
rect 764 979 765 981
rect 761 985 762 987
rect 764 985 765 987
rect 801 359 802 361
rect 804 359 805 361
rect 801 365 802 367
rect 804 365 805 367
rect 381 679 382 681
rect 384 679 385 681
rect 381 685 382 687
rect 384 685 385 687
rect 341 719 342 721
rect 344 719 345 721
rect 341 725 342 727
rect 344 725 345 727
rect 701 919 702 921
rect 704 919 705 921
rect 701 925 702 927
rect 704 925 705 927
rect 741 419 742 421
rect 744 419 745 421
rect 741 425 742 427
rect 744 425 745 427
rect 761 959 762 961
rect 764 959 765 961
rect 761 965 762 967
rect 764 965 765 967
rect 781 779 782 781
rect 784 779 785 781
rect 781 785 782 787
rect 784 785 785 787
rect 901 759 902 761
rect 904 759 905 761
rect 901 765 902 767
rect 904 765 905 767
rect 661 1079 662 1081
rect 664 1079 665 1081
rect 661 1085 662 1087
rect 664 1085 665 1087
rect 601 1019 602 1021
rect 604 1019 605 1021
rect 601 1025 602 1027
rect 604 1025 605 1027
rect 481 559 482 561
rect 484 559 485 561
rect 481 565 482 567
rect 484 565 485 567
rect 541 919 542 921
rect 544 919 545 921
rect 541 925 542 927
rect 544 925 545 927
rect 721 559 722 561
rect 724 559 725 561
rect 721 565 722 567
rect 724 565 725 567
rect 781 479 782 481
rect 784 479 785 481
rect 781 485 782 487
rect 784 485 785 487
rect 941 779 942 781
rect 944 779 945 781
rect 941 785 942 787
rect 944 785 945 787
rect 1001 619 1002 621
rect 1004 619 1005 621
rect 1001 625 1002 627
rect 1004 625 1005 627
rect 621 439 622 441
rect 624 439 625 441
rect 621 445 622 447
rect 624 445 625 447
rect 621 899 622 901
rect 624 899 625 901
rect 621 905 622 907
rect 624 905 625 907
rect 281 719 282 721
rect 284 719 285 721
rect 281 725 282 727
rect 284 725 285 727
rect 921 639 922 641
rect 924 639 925 641
rect 921 645 922 647
rect 924 645 925 647
rect 721 399 722 401
rect 724 399 725 401
rect 721 405 722 407
rect 724 405 725 407
rect 381 799 382 801
rect 384 799 385 801
rect 381 805 382 807
rect 384 805 385 807
rect 861 479 862 481
rect 864 479 865 481
rect 861 485 862 487
rect 864 485 865 487
rect 781 599 782 601
rect 784 599 785 601
rect 781 605 782 607
rect 784 605 785 607
rect 641 579 642 581
rect 644 579 645 581
rect 641 585 642 587
rect 644 585 645 587
rect 341 599 342 601
rect 344 599 345 601
rect 341 605 342 607
rect 344 605 345 607
rect 921 539 922 541
rect 924 539 925 541
rect 921 545 922 547
rect 924 545 925 547
rect 781 379 782 381
rect 784 379 785 381
rect 781 385 782 387
rect 784 385 785 387
rect 521 959 522 961
rect 524 959 525 961
rect 521 965 522 967
rect 524 965 525 967
rect 1021 599 1022 601
rect 1024 599 1025 601
rect 1021 605 1022 607
rect 1024 605 1025 607
rect 721 339 722 341
rect 724 339 725 341
rect 721 345 722 347
rect 724 345 725 347
rect 481 859 482 861
rect 484 859 485 861
rect 481 865 482 867
rect 484 865 485 867
rect 361 679 362 681
rect 364 679 365 681
rect 361 685 362 687
rect 364 685 365 687
rect 301 599 302 601
rect 304 599 305 601
rect 301 605 302 607
rect 304 605 305 607
rect 701 339 702 341
rect 704 339 705 341
rect 701 345 702 347
rect 704 345 705 347
rect 641 979 642 981
rect 644 979 645 981
rect 641 985 642 987
rect 644 985 645 987
rect 361 759 362 761
rect 364 759 365 761
rect 361 765 362 767
rect 364 765 365 767
rect 381 779 382 781
rect 384 779 385 781
rect 381 785 382 787
rect 384 785 385 787
rect 901 679 902 681
rect 904 679 905 681
rect 901 685 902 687
rect 904 685 905 687
rect 781 659 782 661
rect 784 659 785 661
rect 781 665 782 667
rect 784 665 785 667
rect 801 679 802 681
rect 804 679 805 681
rect 801 685 802 687
rect 804 685 805 687
rect 681 719 682 721
rect 684 719 685 721
rect 681 725 682 727
rect 684 725 685 727
rect 501 739 502 741
rect 504 739 505 741
rect 501 745 502 747
rect 504 745 505 747
rect 721 579 722 581
rect 724 579 725 581
rect 721 585 722 587
rect 724 585 725 587
rect 281 699 282 701
rect 284 699 285 701
rect 281 705 282 707
rect 284 705 285 707
rect 841 559 842 561
rect 844 559 845 561
rect 841 565 842 567
rect 844 565 845 567
rect 381 759 382 761
rect 384 759 385 761
rect 381 765 382 767
rect 384 765 385 767
rect 621 639 622 641
rect 624 639 625 641
rect 621 645 622 647
rect 624 645 625 647
rect 541 879 542 881
rect 544 879 545 881
rect 541 885 542 887
rect 544 885 545 887
rect 1021 619 1022 621
rect 1024 619 1025 621
rect 1021 625 1022 627
rect 1024 625 1025 627
rect 781 559 782 561
rect 784 559 785 561
rect 781 565 782 567
rect 784 565 785 567
rect 461 659 462 661
rect 464 659 465 661
rect 461 665 462 667
rect 464 665 465 667
rect 761 539 762 541
rect 764 539 765 541
rect 761 545 762 547
rect 764 545 765 547
rect 421 719 422 721
rect 424 719 425 721
rect 421 725 422 727
rect 424 725 425 727
rect 541 519 542 521
rect 544 519 545 521
rect 541 525 542 527
rect 544 525 545 527
rect 521 819 522 821
rect 524 819 525 821
rect 521 825 522 827
rect 524 825 525 827
rect 961 559 962 561
rect 964 559 965 561
rect 961 565 962 567
rect 964 565 965 567
rect 581 579 582 581
rect 584 579 585 581
rect 581 585 582 587
rect 584 585 585 587
rect 801 759 802 761
rect 804 759 805 761
rect 801 765 802 767
rect 804 765 805 767
rect 881 559 882 561
rect 884 559 885 561
rect 881 565 882 567
rect 884 565 885 567
rect 761 579 762 581
rect 764 579 765 581
rect 761 585 762 587
rect 764 585 765 587
rect 741 839 742 841
rect 744 839 745 841
rect 741 845 742 847
rect 744 845 745 847
rect 641 599 642 601
rect 644 599 645 601
rect 641 605 642 607
rect 644 605 645 607
rect 781 739 782 741
rect 784 739 785 741
rect 781 745 782 747
rect 784 745 785 747
rect 781 719 782 721
rect 784 719 785 721
rect 781 725 782 727
rect 784 725 785 727
rect 601 699 602 701
rect 604 699 605 701
rect 601 705 602 707
rect 604 705 605 707
rect 981 739 982 741
rect 984 739 985 741
rect 981 745 982 747
rect 984 745 985 747
rect 321 799 322 801
rect 324 799 325 801
rect 321 805 322 807
rect 324 805 325 807
rect 901 599 902 601
rect 904 599 905 601
rect 901 605 902 607
rect 904 605 905 607
rect 1001 719 1002 721
rect 1004 719 1005 721
rect 1001 725 1002 727
rect 1004 725 1005 727
rect 581 879 582 881
rect 584 879 585 881
rect 581 885 582 887
rect 584 885 585 887
rect 621 459 622 461
rect 624 459 625 461
rect 621 465 622 467
rect 624 465 625 467
rect 841 439 842 441
rect 844 439 845 441
rect 841 445 842 447
rect 844 445 845 447
rect 801 779 802 781
rect 804 779 805 781
rect 801 785 802 787
rect 804 785 805 787
rect 641 879 642 881
rect 644 879 645 881
rect 641 885 642 887
rect 644 885 645 887
rect 841 919 842 921
rect 844 919 845 921
rect 841 925 842 927
rect 844 925 845 927
rect 701 379 702 381
rect 704 379 705 381
rect 701 385 702 387
rect 704 385 705 387
rect 601 619 602 621
rect 604 619 605 621
rect 601 625 602 627
rect 604 625 605 627
rect 541 659 542 661
rect 544 659 545 661
rect 541 665 542 667
rect 544 665 545 667
rect 641 1059 642 1061
rect 644 1059 645 1061
rect 641 1065 642 1067
rect 644 1065 645 1067
rect 381 819 382 821
rect 384 819 385 821
rect 381 825 382 827
rect 384 825 385 827
rect 621 1079 622 1081
rect 624 1079 625 1081
rect 621 1085 622 1087
rect 624 1085 625 1087
rect 781 959 782 961
rect 784 959 785 961
rect 781 965 782 967
rect 784 965 785 967
rect 661 299 662 301
rect 664 299 665 301
rect 661 305 662 307
rect 664 305 665 307
rect 521 439 522 441
rect 524 439 525 441
rect 521 445 522 447
rect 524 445 525 447
rect 801 439 802 441
rect 804 439 805 441
rect 801 445 802 447
rect 804 445 805 447
rect 341 779 342 781
rect 344 779 345 781
rect 341 785 342 787
rect 344 785 345 787
rect 541 499 542 501
rect 544 499 545 501
rect 541 505 542 507
rect 544 505 545 507
rect 561 699 562 701
rect 564 699 565 701
rect 561 705 562 707
rect 564 705 565 707
rect 441 579 442 581
rect 444 579 445 581
rect 441 585 442 587
rect 444 585 445 587
rect 541 979 542 981
rect 544 979 545 981
rect 541 985 542 987
rect 544 985 545 987
rect 421 619 422 621
rect 424 619 425 621
rect 421 625 422 627
rect 424 625 425 627
rect 301 699 302 701
rect 304 699 305 701
rect 301 705 302 707
rect 304 705 305 707
rect 381 579 382 581
rect 384 579 385 581
rect 381 585 382 587
rect 384 585 385 587
rect 561 999 562 1001
rect 564 999 565 1001
rect 561 1005 562 1007
rect 564 1005 565 1007
rect 661 919 662 921
rect 664 919 665 921
rect 661 925 662 927
rect 664 925 665 927
rect 741 359 742 361
rect 744 359 745 361
rect 741 365 742 367
rect 744 365 745 367
rect 541 579 542 581
rect 544 579 545 581
rect 541 585 542 587
rect 544 585 545 587
rect 421 879 422 881
rect 424 879 425 881
rect 421 885 422 887
rect 424 885 425 887
rect 841 479 842 481
rect 844 479 845 481
rect 841 485 842 487
rect 844 485 845 487
rect 621 499 622 501
rect 624 499 625 501
rect 621 505 622 507
rect 624 505 625 507
rect 601 739 602 741
rect 604 739 605 741
rect 601 745 602 747
rect 604 745 605 747
rect 321 779 322 781
rect 324 779 325 781
rect 321 785 322 787
rect 324 785 325 787
rect 741 979 742 981
rect 744 979 745 981
rect 741 985 742 987
rect 744 985 745 987
rect 881 859 882 861
rect 884 859 885 861
rect 881 865 882 867
rect 884 865 885 867
rect 441 619 442 621
rect 444 619 445 621
rect 441 625 442 627
rect 444 625 445 627
rect 381 559 382 561
rect 384 559 385 561
rect 381 565 382 567
rect 384 565 385 567
rect 561 979 562 981
rect 564 979 565 981
rect 561 985 562 987
rect 564 985 565 987
rect 681 399 682 401
rect 684 399 685 401
rect 681 405 682 407
rect 684 405 685 407
rect 561 399 562 401
rect 564 399 565 401
rect 561 405 562 407
rect 564 405 565 407
rect 621 779 622 781
rect 624 779 625 781
rect 621 785 622 787
rect 624 785 625 787
rect 661 1059 662 1061
rect 664 1059 665 1061
rect 661 1065 662 1067
rect 664 1065 665 1067
rect 861 639 862 641
rect 864 639 865 641
rect 861 645 862 647
rect 864 645 865 647
rect 661 639 662 641
rect 664 639 665 641
rect 661 645 662 647
rect 664 645 665 647
rect 581 379 582 381
rect 584 379 585 381
rect 581 385 582 387
rect 584 385 585 387
rect 601 459 602 461
rect 604 459 605 461
rect 601 465 602 467
rect 604 465 605 467
rect 341 659 342 661
rect 344 659 345 661
rect 341 665 342 667
rect 344 665 345 667
rect 721 1039 722 1041
rect 724 1039 725 1041
rect 721 1045 722 1047
rect 724 1045 725 1047
rect 1041 619 1042 621
rect 1044 619 1045 621
rect 1041 625 1042 627
rect 1044 625 1045 627
rect 821 839 822 841
rect 824 839 825 841
rect 821 845 822 847
rect 824 845 825 847
rect 561 839 562 841
rect 564 839 565 841
rect 561 845 562 847
rect 564 845 565 847
rect 561 459 562 461
rect 564 459 565 461
rect 561 465 562 467
rect 564 465 565 467
rect 901 859 902 861
rect 904 859 905 861
rect 901 865 902 867
rect 904 865 905 867
rect 721 439 722 441
rect 724 439 725 441
rect 721 445 722 447
rect 724 445 725 447
rect 741 879 742 881
rect 744 879 745 881
rect 741 885 742 887
rect 744 885 745 887
rect 701 399 702 401
rect 704 399 705 401
rect 701 405 702 407
rect 704 405 705 407
rect 761 999 762 1001
rect 764 999 765 1001
rect 761 1005 762 1007
rect 764 1005 765 1007
rect 701 459 702 461
rect 704 459 705 461
rect 701 465 702 467
rect 704 465 705 467
rect 481 399 482 401
rect 484 399 485 401
rect 481 405 482 407
rect 484 405 485 407
rect 741 559 742 561
rect 744 559 745 561
rect 741 565 742 567
rect 744 565 745 567
rect 521 859 522 861
rect 524 859 525 861
rect 521 865 522 867
rect 524 865 525 867
rect 901 539 902 541
rect 904 539 905 541
rect 901 545 902 547
rect 904 545 905 547
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
<< labels >>
rlabel pdiffusion 683 703 684 704 0 Cellno = 1
rlabel pdiffusion 583 423 584 424 0 Cellno = 2
rlabel pdiffusion 743 603 744 604 0 Cellno = 3
rlabel pdiffusion 763 523 764 524 0 Cellno = 4
rlabel pdiffusion 643 843 644 844 0 Cellno = 5
rlabel pdiffusion 643 743 644 744 0 Cellno = 6
rlabel pdiffusion 603 923 604 924 0 Cellno = 7
rlabel pdiffusion 503 803 504 804 0 Cellno = 8
rlabel pdiffusion 803 663 804 664 0 Cellno = 9
rlabel pdiffusion 483 643 484 644 0 Cellno = 10
rlabel pdiffusion 843 623 844 624 0 Cellno = 11
rlabel pdiffusion 763 663 764 664 0 Cellno = 12
rlabel pdiffusion 703 703 704 704 0 Cellno = 13
rlabel pdiffusion 523 543 524 544 0 Cellno = 14
rlabel pdiffusion 423 863 424 864 0 Cellno = 15
rlabel pdiffusion 603 903 604 904 0 Cellno = 16
rlabel pdiffusion 443 843 444 844 0 Cellno = 17
rlabel pdiffusion 683 743 684 744 0 Cellno = 18
rlabel pdiffusion 543 543 544 544 0 Cellno = 19
rlabel pdiffusion 863 743 864 744 0 Cellno = 20
rlabel pdiffusion 563 883 564 884 0 Cellno = 21
rlabel pdiffusion 563 603 564 604 0 Cellno = 22
rlabel pdiffusion 643 543 644 544 0 Cellno = 23
rlabel pdiffusion 643 803 644 804 0 Cellno = 24
rlabel pdiffusion 543 803 544 804 0 Cellno = 25
rlabel pdiffusion 583 903 584 904 0 Cellno = 26
rlabel pdiffusion 923 723 924 724 0 Cellno = 27
rlabel pdiffusion 483 763 484 764 0 Cellno = 28
rlabel pdiffusion 683 663 684 664 0 Cellno = 29
rlabel pdiffusion 683 843 684 844 0 Cellno = 30
rlabel pdiffusion 763 483 764 484 0 Cellno = 31
rlabel pdiffusion 403 843 404 844 0 Cellno = 32
rlabel pdiffusion 463 563 464 564 0 Cellno = 33
rlabel pdiffusion 443 723 444 724 0 Cellno = 34
rlabel pdiffusion 603 583 604 584 0 Cellno = 35
rlabel pdiffusion 923 703 924 704 0 Cellno = 36
rlabel pdiffusion 763 623 764 624 0 Cellno = 37
rlabel pdiffusion 703 783 704 784 0 Cellno = 38
rlabel pdiffusion 643 643 644 644 0 Cellno = 39
rlabel pdiffusion 443 703 444 704 0 Cellno = 40
rlabel pdiffusion 603 643 604 644 0 Cellno = 41
rlabel pdiffusion 723 603 724 604 0 Cellno = 42
rlabel pdiffusion 443 903 444 904 0 Cellno = 43
rlabel pdiffusion 603 523 604 524 0 Cellno = 44
rlabel pdiffusion 583 683 584 684 0 Cellno = 45
rlabel pdiffusion 723 683 724 684 0 Cellno = 46
rlabel pdiffusion 803 703 804 704 0 Cellno = 47
rlabel pdiffusion 783 583 784 584 0 Cellno = 48
rlabel pdiffusion 863 603 864 604 0 Cellno = 49
rlabel pdiffusion 503 943 504 944 0 Cellno = 50
rlabel pdiffusion 743 723 744 724 0 Cellno = 51
rlabel pdiffusion 523 763 524 764 0 Cellno = 52
rlabel pdiffusion 843 743 844 744 0 Cellno = 53
rlabel pdiffusion 703 583 704 584 0 Cellno = 54
rlabel pdiffusion 583 543 584 544 0 Cellno = 55
rlabel pdiffusion 783 763 784 764 0 Cellno = 56
rlabel pdiffusion 603 843 604 844 0 Cellno = 57
rlabel pdiffusion 663 443 664 444 0 Cellno = 58
rlabel pdiffusion 783 643 784 644 0 Cellno = 59
rlabel pdiffusion 523 683 524 684 0 Cellno = 60
rlabel pdiffusion 343 683 344 684 0 Cellno = 61
rlabel pdiffusion 483 663 484 664 0 Cellno = 62
rlabel pdiffusion 603 983 604 984 0 Cellno = 63
rlabel pdiffusion 683 603 684 604 0 Cellno = 64
rlabel pdiffusion 683 903 684 904 0 Cellno = 65
rlabel pdiffusion 823 903 824 904 0 Cellno = 66
rlabel pdiffusion 663 783 664 784 0 Cellno = 67
rlabel pdiffusion 683 863 684 864 0 Cellno = 68
rlabel pdiffusion 663 883 664 884 0 Cellno = 69
rlabel pdiffusion 343 703 344 704 0 Cellno = 70
rlabel pdiffusion 543 563 544 564 0 Cellno = 71
rlabel pdiffusion 383 863 384 864 0 Cellno = 72
rlabel pdiffusion 723 743 724 744 0 Cellno = 73
rlabel pdiffusion 523 743 524 744 0 Cellno = 74
rlabel pdiffusion 623 883 624 884 0 Cellno = 75
rlabel pdiffusion 623 383 624 384 0 Cellno = 76
rlabel pdiffusion 663 623 664 624 0 Cellno = 77
rlabel pdiffusion 763 703 764 704 0 Cellno = 78
rlabel pdiffusion 863 503 864 504 0 Cellno = 79
rlabel pdiffusion 503 843 504 844 0 Cellno = 80
rlabel pdiffusion 703 483 704 484 0 Cellno = 81
rlabel pdiffusion 523 563 524 564 0 Cellno = 82
rlabel pdiffusion 963 683 964 684 0 Cellno = 83
rlabel pdiffusion 443 563 444 564 0 Cellno = 84
rlabel pdiffusion 483 783 484 784 0 Cellno = 85
rlabel pdiffusion 483 883 484 884 0 Cellno = 86
rlabel pdiffusion 663 683 664 684 0 Cellno = 87
rlabel pdiffusion 643 463 644 464 0 Cellno = 88
rlabel pdiffusion 843 843 844 844 0 Cellno = 89
rlabel pdiffusion 623 683 624 684 0 Cellno = 90
rlabel pdiffusion 923 783 924 784 0 Cellno = 91
rlabel pdiffusion 443 643 444 644 0 Cellno = 92
rlabel pdiffusion 923 803 924 804 0 Cellno = 93
rlabel pdiffusion 383 603 384 604 0 Cellno = 94
rlabel pdiffusion 803 823 804 824 0 Cellno = 95
rlabel pdiffusion 463 923 464 924 0 Cellno = 96
rlabel pdiffusion 363 543 364 544 0 Cellno = 97
rlabel pdiffusion 663 563 664 564 0 Cellno = 98
rlabel pdiffusion 643 483 644 484 0 Cellno = 99
rlabel pdiffusion 743 623 744 624 0 Cellno = 100
rlabel pdiffusion 663 903 664 904 0 Cellno = 101
rlabel pdiffusion 803 483 804 484 0 Cellno = 102
rlabel pdiffusion 803 723 804 724 0 Cellno = 103
rlabel pdiffusion 463 623 464 624 0 Cellno = 104
rlabel pdiffusion 563 543 564 544 0 Cellno = 105
rlabel pdiffusion 623 723 624 724 0 Cellno = 106
rlabel pdiffusion 803 803 804 804 0 Cellno = 107
rlabel pdiffusion 603 603 604 604 0 Cellno = 108
rlabel pdiffusion 923 843 924 844 0 Cellno = 109
rlabel pdiffusion 483 543 484 544 0 Cellno = 110
rlabel pdiffusion 923 563 924 564 0 Cellno = 111
rlabel pdiffusion 643 703 644 704 0 Cellno = 112
rlabel pdiffusion 643 523 644 524 0 Cellno = 113
rlabel pdiffusion 923 683 924 684 0 Cellno = 114
rlabel pdiffusion 623 763 624 764 0 Cellno = 115
rlabel pdiffusion 423 743 424 744 0 Cellno = 116
rlabel pdiffusion 803 523 804 524 0 Cellno = 117
rlabel pdiffusion 723 463 724 464 0 Cellno = 118
rlabel pdiffusion 923 583 924 584 0 Cellno = 119
rlabel pdiffusion 563 783 564 784 0 Cellno = 120
rlabel pdiffusion 503 383 504 384 0 Cellno = 121
rlabel pdiffusion 943 603 944 604 0 Cellno = 122
rlabel pdiffusion 423 543 424 544 0 Cellno = 123
rlabel pdiffusion 943 623 944 624 0 Cellno = 124
rlabel pdiffusion 563 723 564 724 0 Cellno = 125
rlabel pdiffusion 463 863 464 864 0 Cellno = 126
rlabel pdiffusion 563 823 564 824 0 Cellno = 127
rlabel pdiffusion 743 643 744 644 0 Cellno = 128
rlabel pdiffusion 763 883 764 884 0 Cellno = 129
rlabel pdiffusion 483 683 484 684 0 Cellno = 130
rlabel pdiffusion 843 943 844 944 0 Cellno = 131
rlabel pdiffusion 863 463 864 464 0 Cellno = 132
rlabel pdiffusion 663 603 664 604 0 Cellno = 133
rlabel pdiffusion 483 483 484 484 0 Cellno = 134
rlabel pdiffusion 723 523 724 524 0 Cellno = 135
rlabel pdiffusion 503 583 504 584 0 Cellno = 136
rlabel pdiffusion 363 843 364 844 0 Cellno = 137
rlabel pdiffusion 363 823 364 824 0 Cellno = 138
rlabel pdiffusion 743 523 744 524 0 Cellno = 139
rlabel pdiffusion 843 783 844 784 0 Cellno = 140
rlabel pdiffusion 383 623 384 624 0 Cellno = 141
rlabel pdiffusion 483 843 484 844 0 Cellno = 142
rlabel pdiffusion 563 483 564 484 0 Cellno = 143
rlabel pdiffusion 443 683 444 684 0 Cellno = 144
rlabel pdiffusion 503 703 504 704 0 Cellno = 145
rlabel pdiffusion 523 843 524 844 0 Cellno = 146
rlabel pdiffusion 543 643 544 644 0 Cellno = 147
rlabel pdiffusion 803 563 804 564 0 Cellno = 148
rlabel pdiffusion 563 523 564 524 0 Cellno = 149
rlabel pdiffusion 583 703 584 704 0 Cellno = 150
rlabel pdiffusion 603 803 604 804 0 Cellno = 151
rlabel pdiffusion 823 883 824 884 0 Cellno = 152
rlabel pdiffusion 763 783 764 784 0 Cellno = 153
rlabel pdiffusion 623 963 624 964 0 Cellno = 154
rlabel pdiffusion 483 703 484 704 0 Cellno = 155
rlabel pdiffusion 503 443 504 444 0 Cellno = 156
rlabel pdiffusion 523 643 524 644 0 Cellno = 157
rlabel pdiffusion 763 683 764 684 0 Cellno = 158
rlabel pdiffusion 543 823 544 824 0 Cellno = 159
rlabel pdiffusion 563 383 564 384 0 Cellno = 160
rlabel pdiffusion 863 783 864 784 0 Cellno = 161
rlabel pdiffusion 663 463 664 464 0 Cellno = 162
rlabel pdiffusion 683 303 684 304 0 Cellno = 163
rlabel pdiffusion 643 623 644 624 0 Cellno = 164
rlabel pdiffusion 563 663 564 664 0 Cellno = 165
rlabel pdiffusion 363 603 364 604 0 Cellno = 166
rlabel pdiffusion 643 1023 644 1024 0 Cellno = 167
rlabel pdiffusion 723 823 724 824 0 Cellno = 168
rlabel pdiffusion 763 723 764 724 0 Cellno = 169
rlabel pdiffusion 663 803 664 804 0 Cellno = 170
rlabel pdiffusion 563 683 564 684 0 Cellno = 171
rlabel pdiffusion 463 743 464 744 0 Cellno = 172
rlabel pdiffusion 743 323 744 324 0 Cellno = 173
rlabel pdiffusion 703 523 704 524 0 Cellno = 174
rlabel pdiffusion 503 723 504 724 0 Cellno = 175
rlabel pdiffusion 703 903 704 904 0 Cellno = 176
rlabel pdiffusion 963 583 964 584 0 Cellno = 177
rlabel pdiffusion 743 963 744 964 0 Cellno = 178
rlabel pdiffusion 603 1043 604 1044 0 Cellno = 179
rlabel pdiffusion 763 943 764 944 0 Cellno = 180
rlabel pdiffusion 803 643 804 644 0 Cellno = 181
rlabel pdiffusion 323 763 324 764 0 Cellno = 182
rlabel pdiffusion 823 603 824 604 0 Cellno = 183
rlabel pdiffusion 723 303 724 304 0 Cellno = 184
rlabel pdiffusion 683 463 684 464 0 Cellno = 185
rlabel pdiffusion 823 563 824 564 0 Cellno = 186
rlabel pdiffusion 723 803 724 804 0 Cellno = 187
rlabel pdiffusion 623 923 624 924 0 Cellno = 188
rlabel pdiffusion 363 803 364 804 0 Cellno = 189
rlabel pdiffusion 543 763 544 764 0 Cellno = 190
rlabel pdiffusion 483 503 484 504 0 Cellno = 191
rlabel pdiffusion 623 563 624 564 0 Cellno = 192
rlabel pdiffusion 703 1023 704 1024 0 Cellno = 193
rlabel pdiffusion 863 923 864 924 0 Cellno = 194
rlabel pdiffusion 863 763 864 764 0 Cellno = 195
rlabel pdiffusion 983 683 984 684 0 Cellno = 196
rlabel pdiffusion 423 843 424 844 0 Cellno = 197
rlabel pdiffusion 783 843 784 844 0 Cellno = 198
rlabel pdiffusion 843 463 844 464 0 Cellno = 199
rlabel pdiffusion 503 783 504 784 0 Cellno = 200
rlabel pdiffusion 583 603 584 604 0 Cellno = 201
rlabel pdiffusion 703 323 704 324 0 Cellno = 202
rlabel pdiffusion 563 363 564 364 0 Cellno = 203
rlabel pdiffusion 783 903 784 904 0 Cellno = 204
rlabel pdiffusion 483 443 484 444 0 Cellno = 205
rlabel pdiffusion 803 543 804 544 0 Cellno = 206
rlabel pdiffusion 763 363 764 364 0 Cellno = 207
rlabel pdiffusion 623 483 624 484 0 Cellno = 208
rlabel pdiffusion 843 683 844 684 0 Cellno = 209
rlabel pdiffusion 563 743 564 744 0 Cellno = 210
rlabel pdiffusion 903 623 904 624 0 Cellno = 211
rlabel pdiffusion 443 483 444 484 0 Cellno = 212
rlabel pdiffusion 763 403 764 404 0 Cellno = 213
rlabel pdiffusion 543 723 544 724 0 Cellno = 214
rlabel pdiffusion 663 823 664 824 0 Cellno = 215
rlabel pdiffusion 403 643 404 644 0 Cellno = 216
rlabel pdiffusion 743 1023 744 1024 0 Cellno = 217
rlabel pdiffusion 543 1003 544 1004 0 Cellno = 218
rlabel pdiffusion 783 403 784 404 0 Cellno = 219
rlabel pdiffusion 663 1043 664 1044 0 Cellno = 220
rlabel pdiffusion 603 1063 604 1064 0 Cellno = 221
rlabel pdiffusion 483 743 484 744 0 Cellno = 222
rlabel pdiffusion 463 643 464 644 0 Cellno = 223
rlabel pdiffusion 463 903 464 904 0 Cellno = 224
rlabel pdiffusion 583 463 584 464 0 Cellno = 225
rlabel pdiffusion 643 403 644 404 0 Cellno = 226
rlabel pdiffusion 963 763 964 764 0 Cellno = 227
rlabel pdiffusion 563 963 564 964 0 Cellno = 228
rlabel pdiffusion 683 263 684 264 0 Cellno = 229
rlabel pdiffusion 563 583 564 584 0 Cellno = 230
rlabel pdiffusion 683 923 684 924 0 Cellno = 231
rlabel pdiffusion 503 963 504 964 0 Cellno = 232
rlabel pdiffusion 623 323 624 324 0 Cellno = 233
rlabel pdiffusion 603 383 604 384 0 Cellno = 234
rlabel pdiffusion 883 483 884 484 0 Cellno = 235
rlabel pdiffusion 1003 783 1004 784 0 Cellno = 236
rlabel pdiffusion 263 723 264 724 0 Cellno = 237
rlabel pdiffusion 563 423 564 424 0 Cellno = 238
rlabel pdiffusion 263 743 264 744 0 Cellno = 239
rlabel pdiffusion 863 843 864 844 0 Cellno = 240
rlabel pdiffusion 463 723 464 724 0 Cellno = 241
rlabel pdiffusion 643 723 644 724 0 Cellno = 242
rlabel pdiffusion 723 363 724 364 0 Cellno = 243
rlabel pdiffusion 803 463 804 464 0 Cellno = 244
rlabel pdiffusion 783 883 784 884 0 Cellno = 245
rlabel pdiffusion 903 883 904 884 0 Cellno = 246
rlabel pdiffusion 783 463 784 464 0 Cellno = 247
rlabel pdiffusion 623 1043 624 1044 0 Cellno = 248
rlabel pdiffusion 683 683 684 684 0 Cellno = 249
rlabel pdiffusion 783 543 784 544 0 Cellno = 250
rlabel pdiffusion 703 963 704 964 0 Cellno = 251
rlabel pdiffusion 623 983 624 984 0 Cellno = 252
rlabel pdiffusion 723 643 724 644 0 Cellno = 253
rlabel pdiffusion 703 743 704 744 0 Cellno = 254
rlabel pdiffusion 583 1023 584 1024 0 Cellno = 255
rlabel pdiffusion 263 643 264 644 0 Cellno = 256
rlabel pdiffusion 503 923 504 924 0 Cellno = 257
rlabel pdiffusion 743 463 744 464 0 Cellno = 258
rlabel pdiffusion 283 743 284 744 0 Cellno = 259
rlabel pdiffusion 343 803 344 804 0 Cellno = 260
rlabel pdiffusion 623 403 624 404 0 Cellno = 261
rlabel pdiffusion 783 443 784 444 0 Cellno = 262
rlabel pdiffusion 363 643 364 644 0 Cellno = 263
rlabel pdiffusion 403 663 404 664 0 Cellno = 264
rlabel pdiffusion 523 923 524 924 0 Cellno = 265
rlabel pdiffusion 723 663 724 664 0 Cellno = 266
rlabel pdiffusion 983 763 984 764 0 Cellno = 267
rlabel pdiffusion 903 843 904 844 0 Cellno = 268
rlabel pdiffusion 603 343 604 344 0 Cellno = 269
rlabel pdiffusion 983 563 984 564 0 Cellno = 270
rlabel pdiffusion 683 643 684 644 0 Cellno = 271
rlabel pdiffusion 363 583 364 584 0 Cellno = 272
rlabel pdiffusion 603 683 604 684 0 Cellno = 273
rlabel pdiffusion 923 863 924 864 0 Cellno = 274
rlabel pdiffusion 323 703 324 704 0 Cellno = 275
rlabel pdiffusion 583 783 584 784 0 Cellno = 276
rlabel pdiffusion 703 683 704 684 0 Cellno = 277
rlabel pdiffusion 723 963 724 964 0 Cellno = 278
rlabel pdiffusion 343 743 344 744 0 Cellno = 279
rlabel pdiffusion 603 483 604 484 0 Cellno = 280
rlabel pdiffusion 563 343 564 344 0 Cellno = 281
rlabel pdiffusion 703 803 704 804 0 Cellno = 282
rlabel pdiffusion 943 583 944 584 0 Cellno = 283
rlabel pdiffusion 483 463 484 464 0 Cellno = 284
rlabel pdiffusion 423 483 424 484 0 Cellno = 285
rlabel pdiffusion 483 523 484 524 0 Cellno = 286
rlabel pdiffusion 643 283 644 284 0 Cellno = 287
rlabel pdiffusion 883 603 884 604 0 Cellno = 288
rlabel pdiffusion 643 823 644 824 0 Cellno = 289
rlabel pdiffusion 723 723 724 724 0 Cellno = 290
rlabel pdiffusion 383 543 384 544 0 Cellno = 291
rlabel pdiffusion 443 603 444 604 0 Cellno = 292
rlabel pdiffusion 763 503 764 504 0 Cellno = 293
rlabel pdiffusion 603 423 604 424 0 Cellno = 294
rlabel pdiffusion 623 583 624 584 0 Cellno = 295
rlabel pdiffusion 703 363 704 364 0 Cellno = 296
rlabel pdiffusion 943 543 944 544 0 Cellno = 297
rlabel pdiffusion 343 763 344 764 0 Cellno = 298
rlabel pdiffusion 583 803 584 804 0 Cellno = 299
rlabel pdiffusion 503 663 504 664 0 Cellno = 300
rlabel pdiffusion 503 523 504 524 0 Cellno = 301
rlabel pdiffusion 663 323 664 324 0 Cellno = 302
rlabel pdiffusion 503 603 504 604 0 Cellno = 303
rlabel pdiffusion 663 423 664 424 0 Cellno = 304
rlabel pdiffusion 623 1063 624 1064 0 Cellno = 305
rlabel pdiffusion 523 523 524 524 0 Cellno = 306
rlabel pdiffusion 483 803 484 804 0 Cellno = 307
rlabel pdiffusion 463 543 464 544 0 Cellno = 308
rlabel pdiffusion 723 943 724 944 0 Cellno = 309
rlabel pdiffusion 903 583 904 584 0 Cellno = 310
rlabel pdiffusion 303 663 304 664 0 Cellno = 311
rlabel pdiffusion 523 423 524 424 0 Cellno = 312
rlabel pdiffusion 683 983 684 984 0 Cellno = 313
rlabel pdiffusion 423 683 424 684 0 Cellno = 314
rlabel pdiffusion 623 843 624 844 0 Cellno = 315
rlabel pdiffusion 983 703 984 704 0 Cellno = 316
rlabel pdiffusion 323 623 324 624 0 Cellno = 317
rlabel pdiffusion 383 643 384 644 0 Cellno = 318
rlabel pdiffusion 743 543 744 544 0 Cellno = 319
rlabel pdiffusion 403 623 404 624 0 Cellno = 320
rlabel pdiffusion 583 643 584 644 0 Cellno = 321
rlabel pdiffusion 623 1023 624 1024 0 Cellno = 322
rlabel pdiffusion 723 483 724 484 0 Cellno = 323
rlabel pdiffusion 343 583 344 584 0 Cellno = 324
rlabel pdiffusion 883 643 884 644 0 Cellno = 325
rlabel pdiffusion 583 403 584 404 0 Cellno = 326
rlabel pdiffusion 823 703 824 704 0 Cellno = 327
rlabel pdiffusion 503 763 504 764 0 Cellno = 328
rlabel pdiffusion 443 883 444 884 0 Cellno = 329
rlabel pdiffusion 763 443 764 444 0 Cellno = 330
rlabel pdiffusion 603 303 604 304 0 Cellno = 331
rlabel pdiffusion 963 703 964 704 0 Cellno = 332
rlabel pdiffusion 543 703 544 704 0 Cellno = 333
rlabel pdiffusion 843 903 844 904 0 Cellno = 334
rlabel pdiffusion 563 863 564 864 0 Cellno = 335
rlabel pdiffusion 683 443 684 444 0 Cellno = 336
rlabel pdiffusion 803 883 804 884 0 Cellno = 337
rlabel pdiffusion 783 523 784 524 0 Cellno = 338
rlabel pdiffusion 403 763 404 764 0 Cellno = 339
rlabel pdiffusion 723 283 724 284 0 Cellno = 340
rlabel pdiffusion 503 623 504 624 0 Cellno = 341
rlabel pdiffusion 463 503 464 504 0 Cellno = 342
rlabel pdiffusion 843 723 844 724 0 Cellno = 343
rlabel pdiffusion 623 1003 624 1004 0 Cellno = 344
rlabel pdiffusion 663 1003 664 1004 0 Cellno = 345
rlabel pdiffusion 563 643 564 644 0 Cellno = 346
rlabel pdiffusion 263 603 264 604 0 Cellno = 347
rlabel pdiffusion 403 563 404 564 0 Cellno = 348
rlabel pdiffusion 423 663 424 664 0 Cellno = 349
rlabel pdiffusion 263 663 264 664 0 Cellno = 350
rlabel pdiffusion 663 763 664 764 0 Cellno = 351
rlabel pdiffusion 1023 643 1024 644 0 Cellno = 352
rlabel pdiffusion 643 963 644 964 0 Cellno = 353
rlabel pdiffusion 303 763 304 764 0 Cellno = 354
rlabel pdiffusion 663 863 664 864 0 Cellno = 355
rlabel pdiffusion 963 543 964 544 0 Cellno = 356
rlabel pdiffusion 823 783 824 784 0 Cellno = 357
rlabel pdiffusion 843 883 844 884 0 Cellno = 358
rlabel pdiffusion 743 503 744 504 0 Cellno = 359
rlabel pdiffusion 623 423 624 424 0 Cellno = 360
rlabel pdiffusion 883 903 884 904 0 Cellno = 361
rlabel pdiffusion 283 623 284 624 0 Cellno = 362
rlabel pdiffusion 643 343 644 344 0 Cellno = 363
rlabel pdiffusion 543 623 544 624 0 Cellno = 364
rlabel pdiffusion 483 623 484 624 0 Cellno = 365
rlabel pdiffusion 483 423 484 424 0 Cellno = 366
rlabel pdiffusion 243 683 244 684 0 Cellno = 367
rlabel pdiffusion 603 823 604 824 0 Cellno = 368
rlabel pdiffusion 563 623 564 624 0 Cellno = 369
rlabel pdiffusion 903 823 904 824 0 Cellno = 370
rlabel pdiffusion 803 943 804 944 0 Cellno = 371
rlabel pdiffusion 823 483 824 484 0 Cellno = 372
rlabel pdiffusion 1003 703 1004 704 0 Cellno = 373
rlabel pdiffusion 323 683 324 684 0 Cellno = 374
rlabel pdiffusion 743 383 744 384 0 Cellno = 375
rlabel pdiffusion 943 823 944 824 0 Cellno = 376
rlabel pdiffusion 743 1043 744 1044 0 Cellno = 377
rlabel pdiffusion 423 523 424 524 0 Cellno = 378
rlabel pdiffusion 783 943 784 944 0 Cellno = 379
rlabel pdiffusion 903 483 904 484 0 Cellno = 380
rlabel pdiffusion 743 403 744 404 0 Cellno = 381
rlabel pdiffusion 883 763 884 764 0 Cellno = 382
rlabel pdiffusion 703 1003 704 1004 0 Cellno = 383
rlabel pdiffusion 643 563 644 564 0 Cellno = 384
rlabel pdiffusion 603 323 604 324 0 Cellno = 385
rlabel pdiffusion 763 383 764 384 0 Cellno = 386
rlabel pdiffusion 843 503 844 504 0 Cellno = 387
rlabel pdiffusion 943 563 944 564 0 Cellno = 388
rlabel pdiffusion 1063 663 1064 664 0 Cellno = 389
rlabel pdiffusion 603 723 604 724 0 Cellno = 390
rlabel pdiffusion 443 523 444 524 0 Cellno = 391
rlabel pdiffusion 743 763 744 764 0 Cellno = 392
rlabel pdiffusion 343 563 344 564 0 Cellno = 393
rlabel pdiffusion 363 563 364 564 0 Cellno = 394
rlabel pdiffusion 823 403 824 404 0 Cellno = 395
rlabel pdiffusion 643 1083 644 1084 0 Cellno = 396
rlabel pdiffusion 683 523 684 524 0 Cellno = 397
rlabel pdiffusion 763 643 764 644 0 Cellno = 398
rlabel pdiffusion 823 823 824 824 0 Cellno = 399
rlabel pdiffusion 763 423 764 424 0 Cellno = 400
rlabel pdiffusion 503 883 504 884 0 Cellno = 401
rlabel pdiffusion 623 603 624 604 0 Cellno = 402
rlabel pdiffusion 263 703 264 704 0 Cellno = 403
rlabel pdiffusion 803 503 804 504 0 Cellno = 404
rlabel pdiffusion 423 803 424 804 0 Cellno = 405
rlabel pdiffusion 863 443 864 444 0 Cellno = 406
rlabel pdiffusion 763 1043 764 1044 0 Cellno = 407
rlabel pdiffusion 823 923 824 924 0 Cellno = 408
rlabel pdiffusion 683 783 684 784 0 Cellno = 409
rlabel pdiffusion 663 503 664 504 0 Cellno = 410
rlabel pdiffusion 723 983 724 984 0 Cellno = 411
rlabel pdiffusion 583 663 584 664 0 Cellno = 412
rlabel pdiffusion 943 763 944 764 0 Cellno = 413
rlabel pdiffusion 863 543 864 544 0 Cellno = 414
rlabel pdiffusion 1043 643 1044 644 0 Cellno = 415
rlabel pdiffusion 703 823 704 824 0 Cellno = 416
rlabel pdiffusion 823 863 824 864 0 Cellno = 417
rlabel pdiffusion 963 623 964 624 0 Cellno = 418
rlabel pdiffusion 543 383 544 384 0 Cellno = 419
rlabel pdiffusion 703 943 704 944 0 Cellno = 420
rlabel pdiffusion 643 663 644 664 0 Cellno = 421
rlabel pdiffusion 703 883 704 884 0 Cellno = 422
rlabel pdiffusion 663 543 664 544 0 Cellno = 423
rlabel pdiffusion 743 683 744 684 0 Cellno = 424
rlabel pdiffusion 623 343 624 344 0 Cellno = 425
rlabel pdiffusion 883 583 884 584 0 Cellno = 426
rlabel pdiffusion 703 763 704 764 0 Cellno = 427
rlabel pdiffusion 703 723 704 724 0 Cellno = 428
rlabel pdiffusion 603 563 604 564 0 Cellno = 429
rlabel pdiffusion 583 1043 584 1044 0 Cellno = 430
rlabel pdiffusion 723 543 724 544 0 Cellno = 431
rlabel pdiffusion 623 523 624 524 0 Cellno = 432
rlabel pdiffusion 643 783 644 784 0 Cellno = 433
rlabel pdiffusion 523 583 524 584 0 Cellno = 434
rlabel pdiffusion 523 663 524 664 0 Cellno = 435
rlabel pdiffusion 803 863 804 864 0 Cellno = 436
rlabel pdiffusion 323 603 324 604 0 Cellno = 437
rlabel pdiffusion 543 463 544 464 0 Cellno = 438
rlabel pdiffusion 803 903 804 904 0 Cellno = 439
rlabel pdiffusion 603 1003 604 1004 0 Cellno = 440
rlabel pdiffusion 443 863 444 864 0 Cellno = 441
rlabel pdiffusion 723 423 724 424 0 Cellno = 442
rlabel pdiffusion 583 723 584 724 0 Cellno = 443
rlabel pdiffusion 743 663 744 664 0 Cellno = 444
rlabel pdiffusion 823 623 824 624 0 Cellno = 445
rlabel pdiffusion 363 723 364 724 0 Cellno = 446
rlabel pdiffusion 543 943 544 944 0 Cellno = 447
rlabel pdiffusion 543 683 544 684 0 Cellno = 448
rlabel pdiffusion 963 643 964 644 0 Cellno = 449
rlabel pdiffusion 583 843 584 844 0 Cellno = 450
rlabel pdiffusion 723 903 724 904 0 Cellno = 451
rlabel pdiffusion 663 843 664 844 0 Cellno = 452
rlabel pdiffusion 703 303 704 304 0 Cellno = 453
rlabel pdiffusion 443 763 444 764 0 Cellno = 454
rlabel pdiffusion 443 543 444 544 0 Cellno = 455
rlabel pdiffusion 463 463 464 464 0 Cellno = 456
rlabel pdiffusion 403 703 404 704 0 Cellno = 457
rlabel pdiffusion 683 483 684 484 0 Cellno = 458
rlabel pdiffusion 683 343 684 344 0 Cellno = 459
rlabel pdiffusion 723 923 724 924 0 Cellno = 460
rlabel pdiffusion 543 863 544 864 0 Cellno = 461
rlabel pdiffusion 703 1043 704 1044 0 Cellno = 462
rlabel pdiffusion 783 983 784 984 0 Cellno = 463
rlabel pdiffusion 923 523 924 524 0 Cellno = 464
rlabel pdiffusion 463 603 464 604 0 Cellno = 465
rlabel pdiffusion 863 683 864 684 0 Cellno = 466
rlabel pdiffusion 663 743 664 744 0 Cellno = 467
rlabel pdiffusion 483 583 484 584 0 Cellno = 468
rlabel pdiffusion 823 643 824 644 0 Cellno = 469
rlabel pdiffusion 323 743 324 744 0 Cellno = 470
rlabel pdiffusion 643 903 644 904 0 Cellno = 471
rlabel pdiffusion 663 963 664 964 0 Cellno = 472
rlabel pdiffusion 603 543 604 544 0 Cellno = 473
rlabel pdiffusion 443 463 444 464 0 Cellno = 474
rlabel pdiffusion 683 363 684 364 0 Cellno = 475
rlabel pdiffusion 823 663 824 664 0 Cellno = 476
rlabel pdiffusion 743 863 744 864 0 Cellno = 477
rlabel pdiffusion 623 303 624 304 0 Cellno = 478
rlabel pdiffusion 743 583 744 584 0 Cellno = 479
rlabel pdiffusion 843 663 844 664 0 Cellno = 480
rlabel pdiffusion 243 643 244 644 0 Cellno = 481
rlabel pdiffusion 803 603 804 604 0 Cellno = 482
rlabel pdiffusion 743 743 744 744 0 Cellno = 483
rlabel pdiffusion 683 543 684 544 0 Cellno = 484
rlabel pdiffusion 983 723 984 724 0 Cellno = 485
rlabel pdiffusion 1023 743 1024 744 0 Cellno = 486
rlabel pdiffusion 463 423 464 424 0 Cellno = 487
rlabel pdiffusion 503 403 504 404 0 Cellno = 488
rlabel pdiffusion 403 723 404 724 0 Cellno = 489
rlabel pdiffusion 943 843 944 844 0 Cellno = 490
rlabel pdiffusion 723 383 724 384 0 Cellno = 491
rlabel pdiffusion 303 623 304 624 0 Cellno = 492
rlabel pdiffusion 703 423 704 424 0 Cellno = 493
rlabel pdiffusion 523 803 524 804 0 Cellno = 494
rlabel pdiffusion 523 483 524 484 0 Cellno = 495
rlabel pdiffusion 1003 643 1004 644 0 Cellno = 496
rlabel pdiffusion 463 583 464 584 0 Cellno = 497
rlabel pdiffusion 623 703 624 704 0 Cellno = 498
rlabel pdiffusion 923 743 924 744 0 Cellno = 499
rlabel pdiffusion 563 443 564 444 0 Cellno = 500
rlabel pdiffusion 643 1043 644 1044 0 Cellno = 501
rlabel pdiffusion 843 423 844 424 0 Cellno = 502
rlabel pdiffusion 423 823 424 824 0 Cellno = 503
rlabel pdiffusion 843 703 844 704 0 Cellno = 504
rlabel pdiffusion 603 783 604 784 0 Cellno = 505
rlabel pdiffusion 1063 703 1064 704 0 Cellno = 506
rlabel pdiffusion 723 1023 724 1024 0 Cellno = 507
rlabel pdiffusion 663 1023 664 1024 0 Cellno = 508
rlabel pdiffusion 423 763 424 764 0 Cellno = 509
rlabel pdiffusion 403 803 404 804 0 Cellno = 510
rlabel pdiffusion 503 483 504 484 0 Cellno = 511
rlabel pdiffusion 583 743 584 744 0 Cellno = 512
rlabel pdiffusion 723 1003 724 1004 0 Cellno = 513
rlabel pdiffusion 663 523 664 524 0 Cellno = 514
rlabel pdiffusion 803 623 804 624 0 Cellno = 515
rlabel pdiffusion 723 763 724 764 0 Cellno = 516
rlabel pdiffusion 703 503 704 504 0 Cellno = 517
rlabel pdiffusion 523 983 524 984 0 Cellno = 518
rlabel pdiffusion 623 663 624 664 0 Cellno = 519
rlabel pdiffusion 343 543 344 544 0 Cellno = 520
rlabel pdiffusion 603 503 604 504 0 Cellno = 521
rlabel pdiffusion 943 723 944 724 0 Cellno = 522
rlabel pdiffusion 703 843 704 844 0 Cellno = 523
rlabel pdiffusion 923 663 924 664 0 Cellno = 524
rlabel pdiffusion 843 523 844 524 0 Cellno = 525
rlabel pdiffusion 823 763 824 764 0 Cellno = 526
rlabel pdiffusion 883 823 884 824 0 Cellno = 527
rlabel pdiffusion 463 783 464 784 0 Cellno = 528
rlabel pdiffusion 443 443 444 444 0 Cellno = 529
rlabel pdiffusion 523 623 524 624 0 Cellno = 530
rlabel pdiffusion 443 503 444 504 0 Cellno = 531
rlabel pdiffusion 903 803 904 804 0 Cellno = 532
rlabel pdiffusion 763 463 764 464 0 Cellno = 533
rlabel pdiffusion 963 823 964 824 0 Cellno = 534
rlabel pdiffusion 463 763 464 764 0 Cellno = 535
rlabel pdiffusion 923 623 924 624 0 Cellno = 536
rlabel pdiffusion 483 923 484 924 0 Cellno = 537
rlabel pdiffusion 643 943 644 944 0 Cellno = 538
rlabel pdiffusion 883 703 884 704 0 Cellno = 539
rlabel pdiffusion 603 763 604 764 0 Cellno = 540
rlabel pdiffusion 363 703 364 704 0 Cellno = 541
rlabel pdiffusion 783 503 784 504 0 Cellno = 542
rlabel pdiffusion 283 663 284 664 0 Cellno = 543
rlabel pdiffusion 363 743 364 744 0 Cellno = 544
rlabel pdiffusion 523 783 524 784 0 Cellno = 545
rlabel pdiffusion 403 483 404 484 0 Cellno = 546
rlabel pdiffusion 543 783 544 784 0 Cellno = 547
rlabel pdiffusion 403 743 404 744 0 Cellno = 548
rlabel pdiffusion 563 943 564 944 0 Cellno = 549
rlabel pdiffusion 863 823 864 824 0 Cellno = 550
rlabel pdiffusion 683 623 684 624 0 Cellno = 551
rlabel pdiffusion 903 723 904 724 0 Cellno = 552
rlabel pdiffusion 783 923 784 924 0 Cellno = 553
rlabel pdiffusion 743 943 744 944 0 Cellno = 554
rlabel pdiffusion 1003 663 1004 664 0 Cellno = 555
rlabel pdiffusion 763 343 764 344 0 Cellno = 556
rlabel pdiffusion 683 323 684 324 0 Cellno = 557
rlabel pdiffusion 623 543 624 544 0 Cellno = 558
rlabel pdiffusion 503 563 504 564 0 Cellno = 559
rlabel pdiffusion 963 743 964 744 0 Cellno = 560
rlabel pdiffusion 383 843 384 844 0 Cellno = 561
rlabel pdiffusion 663 583 664 584 0 Cellno = 562
rlabel pdiffusion 623 743 624 744 0 Cellno = 563
rlabel pdiffusion 703 663 704 664 0 Cellno = 564
rlabel pdiffusion 323 663 324 664 0 Cellno = 565
rlabel pdiffusion 323 723 324 724 0 Cellno = 566
rlabel pdiffusion 1043 683 1044 684 0 Cellno = 567
rlabel pdiffusion 543 903 544 904 0 Cellno = 568
rlabel pdiffusion 883 523 884 524 0 Cellno = 569
rlabel pdiffusion 303 643 304 644 0 Cellno = 570
rlabel pdiffusion 423 783 424 784 0 Cellno = 571
rlabel pdiffusion 643 863 644 864 0 Cellno = 572
rlabel pdiffusion 883 503 884 504 0 Cellno = 573
rlabel pdiffusion 403 823 404 824 0 Cellno = 574
rlabel pdiffusion 843 823 844 824 0 Cellno = 575
rlabel pdiffusion 543 403 544 404 0 Cellno = 576
rlabel pdiffusion 543 423 544 424 0 Cellno = 577
rlabel pdiffusion 843 543 844 544 0 Cellno = 578
rlabel pdiffusion 983 803 984 804 0 Cellno = 579
rlabel pdiffusion 523 403 524 404 0 Cellno = 580
rlabel pdiffusion 863 663 864 664 0 Cellno = 581
rlabel pdiffusion 583 323 584 324 0 Cellno = 582
rlabel pdiffusion 763 563 764 564 0 Cellno = 583
rlabel pdiffusion 903 783 904 784 0 Cellno = 584
rlabel pdiffusion 983 623 984 624 0 Cellno = 585
rlabel pdiffusion 683 563 684 564 0 Cellno = 586
rlabel pdiffusion 883 463 884 464 0 Cellno = 587
rlabel pdiffusion 763 843 764 844 0 Cellno = 588
rlabel pdiffusion 923 603 924 604 0 Cellno = 589
rlabel pdiffusion 883 623 884 624 0 Cellno = 590
rlabel pdiffusion 303 743 304 744 0 Cellno = 591
rlabel pdiffusion 1023 663 1024 664 0 Cellno = 592
rlabel pdiffusion 663 983 664 984 0 Cellno = 593
rlabel pdiffusion 803 423 804 424 0 Cellno = 594
rlabel pdiffusion 1003 603 1004 604 0 Cellno = 595
rlabel pdiffusion 863 563 864 564 0 Cellno = 596
rlabel pdiffusion 383 703 384 704 0 Cellno = 597
rlabel pdiffusion 663 663 664 664 0 Cellno = 598
rlabel pdiffusion 523 943 524 944 0 Cellno = 599
rlabel pdiffusion 743 803 744 804 0 Cellno = 600
rlabel pdiffusion 523 503 524 504 0 Cellno = 601
rlabel pdiffusion 543 483 544 484 0 Cellno = 602
rlabel pdiffusion 403 583 404 584 0 Cellno = 603
rlabel pdiffusion 983 643 984 644 0 Cellno = 604
rlabel pdiffusion 463 823 464 824 0 Cellno = 605
rlabel pdiffusion 583 483 584 484 0 Cellno = 606
rlabel pdiffusion 423 583 424 584 0 Cellno = 607
rlabel pdiffusion 403 783 404 784 0 Cellno = 608
rlabel pdiffusion 303 803 304 804 0 Cellno = 609
rlabel pdiffusion 943 523 944 524 0 Cellno = 610
rlabel pdiffusion 583 1003 584 1004 0 Cellno = 611
rlabel pdiffusion 683 283 684 284 0 Cellno = 612
rlabel pdiffusion 883 443 884 444 0 Cellno = 613
rlabel pdiffusion 403 603 404 604 0 Cellno = 614
rlabel pdiffusion 903 563 904 564 0 Cellno = 615
rlabel pdiffusion 1003 763 1004 764 0 Cellno = 616
rlabel pdiffusion 323 643 324 644 0 Cellno = 617
rlabel pdiffusion 683 883 684 884 0 Cellno = 618
rlabel pdiffusion 863 803 864 804 0 Cellno = 619
rlabel pdiffusion 863 703 864 704 0 Cellno = 620
rlabel pdiffusion 1003 683 1004 684 0 Cellno = 621
rlabel pdiffusion 743 703 744 704 0 Cellno = 622
rlabel pdiffusion 303 683 304 684 0 Cellno = 623
rlabel pdiffusion 683 763 684 764 0 Cellno = 624
rlabel pdiffusion 663 403 664 404 0 Cellno = 625
rlabel pdiffusion 383 723 384 724 0 Cellno = 626
rlabel pdiffusion 303 723 304 724 0 Cellno = 627
rlabel pdiffusion 703 983 704 984 0 Cellno = 628
rlabel pdiffusion 543 743 544 744 0 Cellno = 629
rlabel pdiffusion 823 723 824 724 0 Cellno = 630
rlabel pdiffusion 643 763 644 764 0 Cellno = 631
rlabel pdiffusion 763 603 764 604 0 Cellno = 632
rlabel pdiffusion 843 583 844 584 0 Cellno = 633
rlabel pdiffusion 423 603 424 604 0 Cellno = 634
rlabel pdiffusion 743 443 744 444 0 Cellno = 635
rlabel pdiffusion 803 963 804 964 0 Cellno = 636
rlabel pdiffusion 783 863 784 864 0 Cellno = 637
rlabel pdiffusion 683 1023 684 1024 0 Cellno = 638
rlabel pdiffusion 543 963 544 964 0 Cellno = 639
rlabel pdiffusion 983 603 984 604 0 Cellno = 640
rlabel pdiffusion 803 923 804 924 0 Cellno = 641
rlabel pdiffusion 963 663 964 664 0 Cellno = 642
rlabel pdiffusion 643 1003 644 1004 0 Cellno = 643
rlabel pdiffusion 323 583 324 584 0 Cellno = 644
rlabel pdiffusion 583 343 584 344 0 Cellno = 645
rlabel pdiffusion 583 823 584 824 0 Cellno = 646
rlabel pdiffusion 763 823 764 824 0 Cellno = 647
rlabel pdiffusion 583 863 584 864 0 Cellno = 648
rlabel pdiffusion 703 623 704 624 0 Cellno = 649
rlabel pdiffusion 523 603 524 604 0 Cellno = 650
rlabel pdiffusion 583 923 584 924 0 Cellno = 651
rlabel pdiffusion 883 663 884 664 0 Cellno = 652
rlabel pdiffusion 463 883 464 884 0 Cellno = 653
rlabel pdiffusion 523 903 524 904 0 Cellno = 654
rlabel pdiffusion 883 683 884 684 0 Cellno = 655
rlabel pdiffusion 443 783 444 784 0 Cellno = 656
rlabel pdiffusion 403 863 404 864 0 Cellno = 657
rlabel pdiffusion 683 963 684 964 0 Cellno = 658
rlabel pdiffusion 823 463 824 464 0 Cellno = 659
rlabel pdiffusion 723 503 724 504 0 Cellno = 660
rlabel pdiffusion 503 823 504 824 0 Cellno = 661
rlabel pdiffusion 443 803 444 804 0 Cellno = 662
rlabel pdiffusion 763 743 764 744 0 Cellno = 663
rlabel pdiffusion 903 663 904 664 0 Cellno = 664
rlabel pdiffusion 563 803 564 804 0 Cellno = 665
rlabel pdiffusion 923 823 924 824 0 Cellno = 666
rlabel pdiffusion 383 743 384 744 0 Cellno = 667
rlabel pdiffusion 663 703 664 704 0 Cellno = 668
rlabel pdiffusion 543 843 544 844 0 Cellno = 669
rlabel pdiffusion 303 583 304 584 0 Cellno = 670
rlabel pdiffusion 783 703 784 704 0 Cellno = 671
rlabel pdiffusion 483 903 484 904 0 Cellno = 672
rlabel pdiffusion 743 1003 744 1004 0 Cellno = 673
rlabel pdiffusion 663 483 664 484 0 Cellno = 674
rlabel pdiffusion 483 723 484 724 0 Cellno = 675
rlabel pdiffusion 863 583 864 584 0 Cellno = 676
rlabel pdiffusion 423 503 424 504 0 Cellno = 677
rlabel pdiffusion 503 503 504 504 0 Cellno = 678
rlabel pdiffusion 643 683 644 684 0 Cellno = 679
rlabel pdiffusion 903 743 904 744 0 Cellno = 680
rlabel pdiffusion 603 963 604 964 0 Cellno = 681
rlabel pdiffusion 663 723 664 724 0 Cellno = 682
rlabel pdiffusion 783 803 784 804 0 Cellno = 683
rlabel pdiffusion 843 763 844 764 0 Cellno = 684
rlabel pdiffusion 623 823 624 824 0 Cellno = 685
rlabel pdiffusion 383 663 384 664 0 Cellno = 686
rlabel pdiffusion 723 703 724 704 0 Cellno = 687
rlabel pdiffusion 763 763 764 764 0 Cellno = 688
rlabel pdiffusion 643 443 644 444 0 Cellno = 689
rlabel pdiffusion 823 423 824 424 0 Cellno = 690
rlabel pdiffusion 443 663 444 664 0 Cellno = 691
rlabel pdiffusion 783 623 784 624 0 Cellno = 692
rlabel pdiffusion 283 683 284 684 0 Cellno = 693
rlabel pdiffusion 743 923 744 924 0 Cellno = 694
rlabel pdiffusion 423 563 424 564 0 Cellno = 695
rlabel pdiffusion 463 803 464 804 0 Cellno = 696
rlabel pdiffusion 463 483 464 484 0 Cellno = 697
rlabel pdiffusion 843 643 844 644 0 Cellno = 698
rlabel pdiffusion 363 783 364 784 0 Cellno = 699
rlabel pdiffusion 623 943 624 944 0 Cellno = 700
rlabel pdiffusion 883 743 884 744 0 Cellno = 701
rlabel pdiffusion 823 943 824 944 0 Cellno = 702
rlabel pdiffusion 603 863 604 864 0 Cellno = 703
rlabel pdiffusion 683 823 684 824 0 Cellno = 704
rlabel pdiffusion 823 583 824 584 0 Cellno = 705
rlabel pdiffusion 623 623 624 624 0 Cellno = 706
rlabel pdiffusion 603 883 604 884 0 Cellno = 707
rlabel pdiffusion 383 503 384 504 0 Cellno = 708
rlabel pdiffusion 583 503 584 504 0 Cellno = 709
rlabel pdiffusion 883 803 884 804 0 Cellno = 710
rlabel pdiffusion 583 523 584 524 0 Cellno = 711
rlabel pdiffusion 883 783 884 784 0 Cellno = 712
rlabel pdiffusion 523 383 524 384 0 Cellno = 713
rlabel pdiffusion 883 883 884 884 0 Cellno = 714
rlabel pdiffusion 463 703 464 704 0 Cellno = 715
rlabel pdiffusion 283 643 284 644 0 Cellno = 716
rlabel pdiffusion 703 443 704 444 0 Cellno = 717
rlabel pdiffusion 643 363 644 364 0 Cellno = 718
rlabel pdiffusion 863 723 864 724 0 Cellno = 719
rlabel pdiffusion 963 783 964 784 0 Cellno = 720
rlabel pdiffusion 1023 723 1024 724 0 Cellno = 721
rlabel pdiffusion 883 843 884 844 0 Cellno = 722
rlabel pdiffusion 643 423 644 424 0 Cellno = 723
rlabel pdiffusion 843 603 844 604 0 Cellno = 724
rlabel pdiffusion 563 563 564 564 0 Cellno = 725
rlabel pdiffusion 743 903 744 904 0 Cellno = 726
rlabel pdiffusion 583 963 584 964 0 Cellno = 727
rlabel pdiffusion 503 903 504 904 0 Cellno = 728
rlabel pdiffusion 463 523 464 524 0 Cellno = 729
rlabel pdiffusion 683 583 684 584 0 Cellno = 730
rlabel pdiffusion 943 683 944 684 0 Cellno = 731
rlabel pdiffusion 903 523 904 524 0 Cellno = 732
rlabel pdiffusion 603 403 604 404 0 Cellno = 733
rlabel pdiffusion 583 443 584 444 0 Cellno = 734
rlabel pdiffusion 563 503 564 504 0 Cellno = 735
rlabel pdiffusion 503 863 504 864 0 Cellno = 736
rlabel pdiffusion 483 823 484 824 0 Cellno = 737
rlabel pdiffusion 723 863 724 864 0 Cellno = 738
rlabel pdiffusion 603 443 604 444 0 Cellno = 739
rlabel pdiffusion 823 543 824 544 0 Cellno = 740
rlabel pdiffusion 663 363 664 364 0 Cellno = 741
rlabel pdiffusion 583 763 584 764 0 Cellno = 742
rlabel pdiffusion 603 943 604 944 0 Cellno = 743
rlabel pdiffusion 523 703 524 704 0 Cellno = 744
rlabel pdiffusion 683 503 684 504 0 Cellno = 745
rlabel pdiffusion 783 683 784 684 0 Cellno = 746
rlabel pdiffusion 283 603 284 604 0 Cellno = 747
rlabel pdiffusion 683 943 684 944 0 Cellno = 748
rlabel pdiffusion 263 623 264 624 0 Cellno = 749
rlabel pdiffusion 703 543 704 544 0 Cellno = 750
rlabel pdiffusion 643 503 644 504 0 Cellno = 751
rlabel pdiffusion 903 703 904 704 0 Cellno = 752
rlabel pdiffusion 503 683 504 684 0 Cellno = 753
rlabel pdiffusion 483 943 484 944 0 Cellno = 754
rlabel pdiffusion 663 343 664 344 0 Cellno = 755
rlabel pdiffusion 443 743 444 744 0 Cellno = 756
rlabel pdiffusion 723 843 724 844 0 Cellno = 757
rlabel pdiffusion 703 863 704 864 0 Cellno = 758
rlabel pdiffusion 463 443 464 444 0 Cellno = 759
rlabel pdiffusion 743 343 744 344 0 Cellno = 760
rlabel pdiffusion 463 1043 464 1044 0 Cellno = 761
rlabel pdiffusion 643 303 644 304 0 Cellno = 762
rlabel pdiffusion 1043 663 1044 664 0 Cellno = 763
rlabel pdiffusion 503 423 504 424 0 Cellno = 764
rlabel pdiffusion 683 803 684 804 0 Cellno = 765
rlabel pdiffusion 723 623 724 624 0 Cellno = 766
rlabel pdiffusion 343 623 344 624 0 Cellno = 767
rlabel pdiffusion 423 643 424 644 0 Cellno = 768
rlabel pdiffusion 823 383 824 384 0 Cellno = 769
rlabel pdiffusion 363 523 364 524 0 Cellno = 770
rlabel pdiffusion 443 823 444 824 0 Cellno = 771
rlabel pdiffusion 563 923 564 924 0 Cellno = 772
rlabel pdiffusion 823 743 824 744 0 Cellno = 773
rlabel pdiffusion 923 763 924 764 0 Cellno = 774
rlabel pdiffusion 623 863 624 864 0 Cellno = 775
rlabel pdiffusion 683 383 684 384 0 Cellno = 776
rlabel pdiffusion 703 563 704 564 0 Cellno = 777
rlabel pdiffusion 923 503 924 504 0 Cellno = 778
rlabel pdiffusion 543 443 544 444 0 Cellno = 779
rlabel pdiffusion 503 543 504 544 0 Cellno = 780
rlabel pdiffusion 943 743 944 744 0 Cellno = 781
rlabel pdiffusion 843 863 844 864 0 Cellno = 782
rlabel pdiffusion 823 443 824 444 0 Cellno = 783
rlabel pdiffusion 943 643 944 644 0 Cellno = 784
rlabel pdiffusion 523 463 524 464 0 Cellno = 785
rlabel pdiffusion 1003 743 1004 744 0 Cellno = 786
rlabel pdiffusion 683 1003 684 1004 0 Cellno = 787
rlabel pdiffusion 503 643 504 644 0 Cellno = 788
rlabel pdiffusion 963 723 964 724 0 Cellno = 789
rlabel pdiffusion 703 603 704 604 0 Cellno = 790
rlabel pdiffusion 583 563 584 564 0 Cellno = 791
rlabel pdiffusion 763 903 764 904 0 Cellno = 792
rlabel pdiffusion 763 863 764 864 0 Cellno = 793
rlabel pdiffusion 603 663 604 664 0 Cellno = 794
rlabel pdiffusion 863 623 864 624 0 Cellno = 795
rlabel pdiffusion 903 503 904 504 0 Cellno = 796
rlabel pdiffusion 543 603 544 604 0 Cellno = 797
rlabel pdiffusion 683 423 684 424 0 Cellno = 798
rlabel pdiffusion 323 563 324 564 0 Cellno = 799
rlabel pdiffusion 563 903 564 904 0 Cellno = 800
rlabel pdiffusion 1023 683 1024 684 0 Cellno = 801
rlabel pdiffusion 483 603 484 604 0 Cellno = 802
rlabel pdiffusion 863 523 864 524 0 Cellno = 803
rlabel pdiffusion 743 783 744 784 0 Cellno = 804
rlabel pdiffusion 1043 703 1044 704 0 Cellno = 805
rlabel pdiffusion 883 723 884 724 0 Cellno = 806
rlabel pdiffusion 563 763 564 764 0 Cellno = 807
rlabel pdiffusion 823 503 824 504 0 Cellno = 808
rlabel pdiffusion 643 323 644 324 0 Cellno = 809
rlabel pdiffusion 763 803 764 804 0 Cellno = 810
rlabel pdiffusion 683 1043 684 1044 0 Cellno = 811
rlabel pdiffusion 643 923 644 924 0 Cellno = 812
rlabel pdiffusion 883 543 884 544 0 Cellno = 813
rlabel pdiffusion 623 803 624 804 0 Cellno = 814
rlabel pdiffusion 383 523 384 524 0 Cellno = 815
rlabel pdiffusion 583 623 584 624 0 Cellno = 816
rlabel pdiffusion 963 603 964 604 0 Cellno = 817
rlabel pdiffusion 743 483 744 484 0 Cellno = 818
rlabel pdiffusion 803 583 804 584 0 Cellno = 819
rlabel pdiffusion 423 463 424 464 0 Cellno = 820
rlabel pdiffusion 503 463 504 464 0 Cellno = 821
rlabel pdiffusion 723 783 724 784 0 Cellno = 822
rlabel pdiffusion 583 943 584 944 0 Cellno = 823
rlabel pdiffusion 643 383 644 384 0 Cellno = 824
rlabel pdiffusion 903 643 904 644 0 Cellno = 825
rlabel pdiffusion 783 823 784 824 0 Cellno = 826
rlabel pdiffusion 343 823 344 824 0 Cellno = 827
rlabel pdiffusion 623 283 624 284 0 Cellno = 828
rlabel pdiffusion 583 363 584 364 0 Cellno = 829
rlabel pdiffusion 803 743 804 744 0 Cellno = 830
rlabel pdiffusion 743 823 744 824 0 Cellno = 831
rlabel pdiffusion 243 703 244 704 0 Cellno = 832
rlabel pdiffusion 463 683 464 684 0 Cellno = 833
rlabel pdiffusion 943 703 944 704 0 Cellno = 834
rlabel pdiffusion 763 923 764 924 0 Cellno = 835
rlabel pdiffusion 803 843 804 844 0 Cellno = 836
rlabel pdiffusion 603 363 604 364 0 Cellno = 837
rlabel pdiffusion 823 523 824 524 0 Cellno = 838
rlabel pdiffusion 843 803 844 804 0 Cellno = 839
rlabel pdiffusion 523 723 524 724 0 Cellno = 840
rlabel pdiffusion 363 623 364 624 0 Cellno = 841
rlabel pdiffusion 703 643 704 644 0 Cellno = 842
rlabel pdiffusion 463 843 464 844 0 Cellno = 843
rlabel pdiffusion 363 663 364 664 0 Cellno = 844
rlabel pdiffusion 723 323 724 324 0 Cellno = 845
rlabel pdiffusion 343 643 344 644 0 Cellno = 846
rlabel pdiffusion 403 683 404 684 0 Cellno = 847
rlabel pdiffusion 983 583 984 584 0 Cellno = 848
rlabel pdiffusion 563 1023 564 1024 0 Cellno = 849
rlabel pdiffusion 783 423 784 424 0 Cellno = 850
rlabel pdiffusion 803 403 804 404 0 Cellno = 851
rlabel pdiffusion 663 383 664 384 0 Cellno = 852
rlabel pdiffusion 403 543 404 544 0 Cellno = 853
rlabel pdiffusion 403 523 404 524 0 Cellno = 854
rlabel pdiffusion 423 703 424 704 0 Cellno = 855
rlabel pdiffusion 863 903 864 904 0 Cellno = 856
rlabel pdiffusion 523 883 524 884 0 Cellno = 857
rlabel pdiffusion 823 683 824 684 0 Cellno = 858
rlabel pdiffusion 863 883 864 884 0 Cellno = 859
rlabel pdiffusion 943 803 944 804 0 Cellno = 860
rlabel pdiffusion 583 983 584 984 0 Cellno = 861
rlabel pdiffusion 623 363 624 364 0 Cellno = 862
rlabel pdiffusion 983 663 984 664 0 Cellno = 863
rlabel pdiffusion 863 863 864 864 0 Cellno = 864
rlabel pdiffusion 663 943 664 944 0 Cellno = 865
rlabel pdiffusion 723 883 724 884 0 Cellno = 866
rlabel pdiffusion 823 803 824 804 0 Cellno = 867
rlabel pdiffusion 763 983 764 984 0 Cellno = 868
rlabel pdiffusion 803 363 804 364 0 Cellno = 869
rlabel pdiffusion 383 683 384 684 0 Cellno = 870
rlabel pdiffusion 343 723 344 724 0 Cellno = 871
rlabel pdiffusion 703 923 704 924 0 Cellno = 872
rlabel pdiffusion 743 423 744 424 0 Cellno = 873
rlabel pdiffusion 763 963 764 964 0 Cellno = 874
rlabel pdiffusion 783 783 784 784 0 Cellno = 875
rlabel pdiffusion 903 763 904 764 0 Cellno = 876
rlabel pdiffusion 663 1083 664 1084 0 Cellno = 877
rlabel pdiffusion 603 1023 604 1024 0 Cellno = 878
rlabel pdiffusion 483 563 484 564 0 Cellno = 879
rlabel pdiffusion 543 923 544 924 0 Cellno = 880
rlabel pdiffusion 723 563 724 564 0 Cellno = 881
rlabel pdiffusion 783 483 784 484 0 Cellno = 882
rlabel pdiffusion 943 783 944 784 0 Cellno = 883
rlabel pdiffusion 1003 623 1004 624 0 Cellno = 884
rlabel pdiffusion 623 443 624 444 0 Cellno = 885
rlabel pdiffusion 623 903 624 904 0 Cellno = 886
rlabel pdiffusion 283 723 284 724 0 Cellno = 887
rlabel pdiffusion 923 643 924 644 0 Cellno = 888
rlabel pdiffusion 723 403 724 404 0 Cellno = 889
rlabel pdiffusion 383 803 384 804 0 Cellno = 890
rlabel pdiffusion 863 483 864 484 0 Cellno = 891
rlabel pdiffusion 783 603 784 604 0 Cellno = 892
rlabel pdiffusion 643 583 644 584 0 Cellno = 893
rlabel pdiffusion 343 603 344 604 0 Cellno = 894
rlabel pdiffusion 923 543 924 544 0 Cellno = 895
rlabel pdiffusion 783 383 784 384 0 Cellno = 896
rlabel pdiffusion 523 963 524 964 0 Cellno = 897
rlabel pdiffusion 1023 603 1024 604 0 Cellno = 898
rlabel pdiffusion 723 343 724 344 0 Cellno = 899
rlabel pdiffusion 483 863 484 864 0 Cellno = 900
rlabel pdiffusion 363 683 364 684 0 Cellno = 901
rlabel pdiffusion 303 603 304 604 0 Cellno = 902
rlabel pdiffusion 703 343 704 344 0 Cellno = 903
rlabel pdiffusion 643 983 644 984 0 Cellno = 904
rlabel pdiffusion 363 763 364 764 0 Cellno = 905
rlabel pdiffusion 383 783 384 784 0 Cellno = 906
rlabel pdiffusion 903 683 904 684 0 Cellno = 907
rlabel pdiffusion 783 663 784 664 0 Cellno = 908
rlabel pdiffusion 803 683 804 684 0 Cellno = 909
rlabel pdiffusion 683 723 684 724 0 Cellno = 910
rlabel pdiffusion 503 743 504 744 0 Cellno = 911
rlabel pdiffusion 723 583 724 584 0 Cellno = 912
rlabel pdiffusion 283 703 284 704 0 Cellno = 913
rlabel pdiffusion 843 563 844 564 0 Cellno = 914
rlabel pdiffusion 383 763 384 764 0 Cellno = 915
rlabel pdiffusion 623 643 624 644 0 Cellno = 916
rlabel pdiffusion 543 883 544 884 0 Cellno = 917
rlabel pdiffusion 1023 623 1024 624 0 Cellno = 918
rlabel pdiffusion 783 563 784 564 0 Cellno = 919
rlabel pdiffusion 463 663 464 664 0 Cellno = 920
rlabel pdiffusion 763 543 764 544 0 Cellno = 921
rlabel pdiffusion 423 723 424 724 0 Cellno = 922
rlabel pdiffusion 543 523 544 524 0 Cellno = 923
rlabel pdiffusion 523 823 524 824 0 Cellno = 924
rlabel pdiffusion 963 563 964 564 0 Cellno = 925
rlabel pdiffusion 583 583 584 584 0 Cellno = 926
rlabel pdiffusion 803 763 804 764 0 Cellno = 927
rlabel pdiffusion 883 563 884 564 0 Cellno = 928
rlabel pdiffusion 763 583 764 584 0 Cellno = 929
rlabel pdiffusion 743 843 744 844 0 Cellno = 930
rlabel pdiffusion 643 603 644 604 0 Cellno = 931
rlabel pdiffusion 783 743 784 744 0 Cellno = 932
rlabel pdiffusion 783 723 784 724 0 Cellno = 933
rlabel pdiffusion 603 703 604 704 0 Cellno = 934
rlabel pdiffusion 983 743 984 744 0 Cellno = 935
rlabel pdiffusion 323 803 324 804 0 Cellno = 936
rlabel pdiffusion 903 603 904 604 0 Cellno = 937
rlabel pdiffusion 1003 723 1004 724 0 Cellno = 938
rlabel pdiffusion 583 883 584 884 0 Cellno = 939
rlabel pdiffusion 623 463 624 464 0 Cellno = 940
rlabel pdiffusion 843 443 844 444 0 Cellno = 941
rlabel pdiffusion 803 783 804 784 0 Cellno = 942
rlabel pdiffusion 643 883 644 884 0 Cellno = 943
rlabel pdiffusion 843 923 844 924 0 Cellno = 944
rlabel pdiffusion 703 383 704 384 0 Cellno = 945
rlabel pdiffusion 603 623 604 624 0 Cellno = 946
rlabel pdiffusion 543 663 544 664 0 Cellno = 947
rlabel pdiffusion 643 1063 644 1064 0 Cellno = 948
rlabel pdiffusion 383 823 384 824 0 Cellno = 949
rlabel pdiffusion 623 1083 624 1084 0 Cellno = 950
rlabel pdiffusion 783 963 784 964 0 Cellno = 951
rlabel pdiffusion 663 303 664 304 0 Cellno = 952
rlabel pdiffusion 523 443 524 444 0 Cellno = 953
rlabel pdiffusion 803 443 804 444 0 Cellno = 954
rlabel pdiffusion 343 783 344 784 0 Cellno = 955
rlabel pdiffusion 543 503 544 504 0 Cellno = 956
rlabel pdiffusion 563 703 564 704 0 Cellno = 957
rlabel pdiffusion 443 583 444 584 0 Cellno = 958
rlabel pdiffusion 543 983 544 984 0 Cellno = 959
rlabel pdiffusion 423 623 424 624 0 Cellno = 960
rlabel pdiffusion 303 703 304 704 0 Cellno = 961
rlabel pdiffusion 383 583 384 584 0 Cellno = 962
rlabel pdiffusion 563 1003 564 1004 0 Cellno = 963
rlabel pdiffusion 663 923 664 924 0 Cellno = 964
rlabel pdiffusion 743 363 744 364 0 Cellno = 965
rlabel pdiffusion 543 583 544 584 0 Cellno = 966
rlabel pdiffusion 423 883 424 884 0 Cellno = 967
rlabel pdiffusion 843 483 844 484 0 Cellno = 968
rlabel pdiffusion 623 503 624 504 0 Cellno = 969
rlabel pdiffusion 603 743 604 744 0 Cellno = 970
rlabel pdiffusion 323 783 324 784 0 Cellno = 971
rlabel pdiffusion 743 983 744 984 0 Cellno = 972
rlabel pdiffusion 883 863 884 864 0 Cellno = 973
rlabel pdiffusion 443 623 444 624 0 Cellno = 974
rlabel pdiffusion 383 563 384 564 0 Cellno = 975
rlabel pdiffusion 563 983 564 984 0 Cellno = 976
rlabel pdiffusion 683 403 684 404 0 Cellno = 977
rlabel pdiffusion 563 403 564 404 0 Cellno = 978
rlabel pdiffusion 623 783 624 784 0 Cellno = 979
rlabel pdiffusion 663 1063 664 1064 0 Cellno = 980
rlabel pdiffusion 863 643 864 644 0 Cellno = 981
rlabel pdiffusion 663 643 664 644 0 Cellno = 982
rlabel pdiffusion 583 383 584 384 0 Cellno = 983
rlabel pdiffusion 603 463 604 464 0 Cellno = 984
rlabel pdiffusion 343 663 344 664 0 Cellno = 985
rlabel pdiffusion 723 1043 724 1044 0 Cellno = 986
rlabel pdiffusion 1043 623 1044 624 0 Cellno = 987
rlabel pdiffusion 823 843 824 844 0 Cellno = 988
rlabel pdiffusion 563 843 564 844 0 Cellno = 989
rlabel pdiffusion 563 463 564 464 0 Cellno = 990
rlabel pdiffusion 903 863 904 864 0 Cellno = 991
rlabel pdiffusion 723 443 724 444 0 Cellno = 992
rlabel pdiffusion 743 883 744 884 0 Cellno = 993
rlabel pdiffusion 703 403 704 404 0 Cellno = 994
rlabel pdiffusion 763 1003 764 1004 0 Cellno = 995
rlabel pdiffusion 703 463 704 464 0 Cellno = 996
rlabel pdiffusion 483 403 484 404 0 Cellno = 997
rlabel pdiffusion 743 563 744 564 0 Cellno = 998
rlabel pdiffusion 523 863 524 864 0 Cellno = 999
rlabel pdiffusion 903 543 904 544 0 Cellno = 1000
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1001
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1002
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1003
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1004
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1005
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1006
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1007
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1008
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1009
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1010
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1011
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1012
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1013
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1014
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1015
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1016
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1017
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1018
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1019
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1020
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1021
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1022
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1023
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1024
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1025
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1026
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1027
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1028
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1029
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1030
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1031
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1032
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1033
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1034
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1035
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1036
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1037
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1038
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1039
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1040
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1041
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1042
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1043
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1044
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1045
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1046
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1047
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1048
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1049
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1050
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1051
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1052
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1053
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1054
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1055
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1056
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1057
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1058
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1059
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1060
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1061
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1062
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1063
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1064
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1065
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1066
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1067
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1068
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1069
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1070
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1071
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1072
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1073
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1074
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1075
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1076
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1077
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1078
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1079
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1080
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1081
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1082
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1083
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1084
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1085
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1086
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1087
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1088
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1089
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1090
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1091
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1092
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1093
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1094
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1095
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1096
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1097
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1098
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1099
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1100
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1101
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1102
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1103
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1104
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1105
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1106
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1107
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1108
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1109
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1110
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1111
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1112
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1113
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1114
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1115
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1116
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1117
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1118
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1119
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1120
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1121
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1122
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1123
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1124
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1125
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1126
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1127
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1128
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1129
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1130
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1131
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1132
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1133
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1134
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1135
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1136
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1137
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1138
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1139
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1140
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1141
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1142
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1143
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1144
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1145
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1146
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1147
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1148
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1149
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1150
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1151
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1152
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1153
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1154
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1155
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1156
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1157
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1158
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1159
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1160
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1161
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1162
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1163
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1164
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1165
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1166
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1167
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1168
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1169
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1170
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1171
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1172
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1173
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1174
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1175
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1176
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1177
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1178
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1179
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1180
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1181
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1182
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1183
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1184
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1185
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1186
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1187
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1188
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1189
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1190
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1191
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1192
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1193
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1194
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1195
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1196
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1197
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1198
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1199
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1200
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1201
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1202
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1203
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1204
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1205
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1206
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1207
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1208
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1209
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1210
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1211
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1212
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1213
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1214
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1215
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1216
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1217
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1218
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1219
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1220
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1221
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1222
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1223
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1224
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1225
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1226
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1227
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1228
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1229
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1230
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1231
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1232
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1233
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1234
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1235
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1236
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1237
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1238
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1239
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1240
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1241
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1242
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1243
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1244
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1245
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1246
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1247
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1248
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1249
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1250
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1251
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1252
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1253
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1254
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1255
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1256
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1257
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1258
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1259
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1260
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1261
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1262
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1263
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1264
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1265
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1266
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1267
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1268
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1269
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1270
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1271
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1272
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1273
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1274
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1275
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1276
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1277
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1278
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1279
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1280
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1281
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1282
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1283
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1284
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1285
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1286
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1287
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1288
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1289
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1290
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1291
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1292
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1293
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1294
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1295
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1296
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1297
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1298
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1299
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1300
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1301
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1302
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1303
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1304
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1305
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1306
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1307
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1308
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1309
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1310
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1311
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1312
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1313
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1314
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1315
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1316
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1317
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1318
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1319
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1320
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1321
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1322
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1323
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1324
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1325
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1326
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1327
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1328
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1329
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1330
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1331
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1332
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1333
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1334
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1335
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1336
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1337
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1338
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1339
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1340
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1341
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1342
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1343
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1344
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1345
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1346
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1347
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1348
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1349
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1350
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1351
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1352
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1353
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1354
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1355
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1356
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1357
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1358
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1359
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1360
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1361
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1362
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1363
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1364
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1365
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1366
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1367
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1368
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1369
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1370
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1371
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1372
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1373
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1374
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1375
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1376
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1377
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1378
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1379
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1380
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1381
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1382
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1383
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1384
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1385
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1386
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1387
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1388
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1389
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1390
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1391
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1392
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1393
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1394
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1395
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1396
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1397
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1398
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1399
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1400
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1401
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1402
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1403
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1404
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1405
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1406
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1407
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1408
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1409
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1410
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1411
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1412
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1413
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1414
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1415
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1416
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1417
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1418
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1419
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1420
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1421
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1422
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1423
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1424
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1425
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1426
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1427
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1428
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1429
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1430
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1431
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1432
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1433
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1434
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1435
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1436
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1437
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1438
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1439
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1440
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1441
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1442
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1443
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1444
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1445
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1446
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1447
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1448
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1449
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1450
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1451
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1452
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1453
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1454
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1455
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1456
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1457
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1458
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1459
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1460
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1461
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1462
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1463
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1464
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1465
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1466
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1467
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1468
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1469
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1470
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1471
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1472
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1473
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1474
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1475
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1476
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1477
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1478
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1479
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1480
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1481
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1482
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1483
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1484
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1485
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1486
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1487
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1488
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1489
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1490
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1491
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1492
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1493
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1494
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1495
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1496
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1497
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1498
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1499
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1500
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1501
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1502
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1503
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1504
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1505
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1506
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1507
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1508
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1509
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1510
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1511
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1512
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1513
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1514
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1515
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1516
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1517
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1518
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1519
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1520
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1521
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1522
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1523
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1524
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1525
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1526
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1527
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1528
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1529
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1530
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1531
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1532
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1533
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1534
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1535
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1536
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1537
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1538
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1539
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1540
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1541
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1542
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1543
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1544
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1545
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1546
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1547
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1548
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1549
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1550
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1551
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1552
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1553
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1554
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1555
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1556
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1557
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1558
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1559
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1560
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1561
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1562
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1563
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1564
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1565
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1566
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1567
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1568
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1569
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1570
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1571
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1572
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1573
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1574
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1575
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1576
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1577
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1578
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1579
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1580
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1581
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1582
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1583
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1584
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1585
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1586
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1587
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1588
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1589
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1590
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1591
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1592
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1593
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1594
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1595
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1596
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1597
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1598
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1599
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1600
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1601
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1602
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1603
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1604
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1605
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1606
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1607
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1608
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1609
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1610
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1611
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1612
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1613
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1614
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1615
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1616
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1617
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1618
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1619
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1620
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1621
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1622
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1623
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1624
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1625
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1626
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1627
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1628
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1629
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1630
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1631
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1632
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1633
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1634
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1635
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1636
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1637
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1638
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1639
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1640
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1641
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1642
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1643
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1644
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1645
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1646
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1647
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1648
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1649
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1650
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1651
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1652
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1653
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1654
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1655
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1656
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1657
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1658
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1659
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1660
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1661
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1662
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1663
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1664
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1665
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1666
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1667
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1668
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1669
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1670
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1671
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1672
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1673
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1674
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1675
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1676
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1677
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1678
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1679
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1680
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1681
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1682
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1683
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1684
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1685
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1686
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1687
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1688
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1689
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1690
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1691
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1692
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1693
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1694
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1695
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1696
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1697
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1698
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1699
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1700
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1701
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1702
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1703
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1704
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1705
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1706
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1707
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1708
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1709
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1710
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1711
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1712
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1713
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1714
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1715
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1716
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1717
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1718
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1719
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1720
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1721
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1722
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1723
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1724
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1725
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1726
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1727
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1728
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1729
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1730
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1731
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1732
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1733
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1734
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1735
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1736
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1737
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1738
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1739
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1740
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1741
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1742
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1743
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1744
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1745
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1746
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1747
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1748
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1749
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1750
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1751
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1752
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1753
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1754
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1755
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1756
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1757
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1758
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1759
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1760
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1761
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1762
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1763
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1764
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1765
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1766
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1767
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1768
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1769
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1770
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1771
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1772
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1773
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1774
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1775
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1776
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1777
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1778
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1779
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1780
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1781
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1782
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1783
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1784
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1785
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1786
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1787
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1788
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1789
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1790
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1791
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1792
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1793
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1794
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1795
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1796
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1797
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1798
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1799
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1800
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1801
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1802
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1803
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1804
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1805
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1806
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1807
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1808
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1809
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1810
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1811
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1812
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1813
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1814
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1815
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1816
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1817
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1818
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1819
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1820
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1821
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1822
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1823
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1824
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1825
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1826
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1827
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1828
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1829
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1830
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1831
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1832
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1833
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1834
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1835
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1836
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1837
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1838
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1839
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1840
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1841
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1842
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1843
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1844
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1845
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1846
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1847
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1848
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1849
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1850
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1851
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1852
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1853
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1854
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1855
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1856
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1857
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1858
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1859
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1860
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1861
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1862
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1863
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1864
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1865
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1866
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1867
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1868
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1869
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1870
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1871
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1872
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1873
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1874
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1875
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1876
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1877
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1878
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1879
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1880
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1881
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1882
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1883
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1884
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1885
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1886
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1887
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1888
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1889
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1890
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1891
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1892
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1893
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1894
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1895
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1896
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1897
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1898
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1899
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1900
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1901
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1902
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1903
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1904
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1905
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1906
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1907
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1908
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1909
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1910
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1911
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1912
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1913
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1914
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1915
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1916
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1917
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1918
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1919
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1920
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1921
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1922
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1923
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1924
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1925
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1926
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1927
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1928
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1929
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1930
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1931
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1932
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1933
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1934
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1935
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1936
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1937
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1938
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1939
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1940
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1941
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1942
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1943
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1944
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1945
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1946
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1947
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1948
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1949
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1950
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1951
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1952
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1953
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1954
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1955
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1956
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1957
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1958
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1959
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1960
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1961
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1962
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1963
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1964
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1965
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1966
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1967
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1968
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1969
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1970
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1971
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1972
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1973
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1974
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1975
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1976
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1977
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1978
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1979
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1980
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1981
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1982
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1983
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1984
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1985
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1986
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1987
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1988
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1989
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1990
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1991
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1992
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1993
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1994
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1995
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1996
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1997
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1998
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1999
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 2000
<< end >>
