magic
tech scmos
timestamp
<< pdiffusion >>
rect 360 260 361 261
rect 362 260 363 261
rect 363 260 364 261
rect 365 260 366 261
rect 360 261 366 265
rect 360 265 361 266
rect 362 265 363 266
rect 363 265 364 266
rect 365 265 366 266
rect 720 420 721 421
rect 722 420 723 421
rect 723 420 724 421
rect 725 420 726 421
rect 720 421 726 425
rect 720 425 721 426
rect 722 425 723 426
rect 723 425 724 426
rect 725 425 726 426
rect 200 380 201 381
rect 202 380 203 381
rect 203 380 204 381
rect 205 380 206 381
rect 200 381 206 385
rect 200 385 201 386
rect 202 385 203 386
rect 203 385 204 386
rect 205 385 206 386
rect 740 480 741 481
rect 742 480 743 481
rect 743 480 744 481
rect 745 480 746 481
rect 740 481 746 485
rect 740 485 741 486
rect 742 485 743 486
rect 743 485 744 486
rect 745 485 746 486
rect 620 820 621 821
rect 622 820 623 821
rect 623 820 624 821
rect 625 820 626 821
rect 620 821 626 825
rect 620 825 621 826
rect 622 825 623 826
rect 623 825 624 826
rect 625 825 626 826
rect 260 540 261 541
rect 262 540 263 541
rect 263 540 264 541
rect 265 540 266 541
rect 260 541 266 545
rect 260 545 261 546
rect 262 545 263 546
rect 263 545 264 546
rect 265 545 266 546
rect 380 400 381 401
rect 382 400 383 401
rect 383 400 384 401
rect 385 400 386 401
rect 380 401 386 405
rect 380 405 381 406
rect 382 405 383 406
rect 383 405 384 406
rect 385 405 386 406
rect 500 420 501 421
rect 502 420 503 421
rect 503 420 504 421
rect 505 420 506 421
rect 500 421 506 425
rect 500 425 501 426
rect 502 425 503 426
rect 503 425 504 426
rect 505 425 506 426
rect 260 360 261 361
rect 262 360 263 361
rect 263 360 264 361
rect 265 360 266 361
rect 260 361 266 365
rect 260 365 261 366
rect 262 365 263 366
rect 263 365 264 366
rect 265 365 266 366
rect 260 660 261 661
rect 262 660 263 661
rect 263 660 264 661
rect 265 660 266 661
rect 260 661 266 665
rect 260 665 261 666
rect 262 665 263 666
rect 263 665 264 666
rect 265 665 266 666
rect 760 660 761 661
rect 762 660 763 661
rect 763 660 764 661
rect 765 660 766 661
rect 760 661 766 665
rect 760 665 761 666
rect 762 665 763 666
rect 763 665 764 666
rect 765 665 766 666
rect 380 660 381 661
rect 382 660 383 661
rect 383 660 384 661
rect 385 660 386 661
rect 380 661 386 665
rect 380 665 381 666
rect 382 665 383 666
rect 383 665 384 666
rect 385 665 386 666
rect 480 800 481 801
rect 482 800 483 801
rect 483 800 484 801
rect 485 800 486 801
rect 480 801 486 805
rect 480 805 481 806
rect 482 805 483 806
rect 483 805 484 806
rect 485 805 486 806
rect 740 680 741 681
rect 742 680 743 681
rect 743 680 744 681
rect 745 680 746 681
rect 740 681 746 685
rect 740 685 741 686
rect 742 685 743 686
rect 743 685 744 686
rect 745 685 746 686
rect 180 480 181 481
rect 182 480 183 481
rect 183 480 184 481
rect 185 480 186 481
rect 180 481 186 485
rect 180 485 181 486
rect 182 485 183 486
rect 183 485 184 486
rect 185 485 186 486
rect 600 620 601 621
rect 602 620 603 621
rect 603 620 604 621
rect 605 620 606 621
rect 600 621 606 625
rect 600 625 601 626
rect 602 625 603 626
rect 603 625 604 626
rect 605 625 606 626
rect 860 540 861 541
rect 862 540 863 541
rect 863 540 864 541
rect 865 540 866 541
rect 860 541 866 545
rect 860 545 861 546
rect 862 545 863 546
rect 863 545 864 546
rect 865 545 866 546
rect 560 580 561 581
rect 562 580 563 581
rect 563 580 564 581
rect 565 580 566 581
rect 560 581 566 585
rect 560 585 561 586
rect 562 585 563 586
rect 563 585 564 586
rect 565 585 566 586
rect 660 620 661 621
rect 662 620 663 621
rect 663 620 664 621
rect 665 620 666 621
rect 660 621 666 625
rect 660 625 661 626
rect 662 625 663 626
rect 663 625 664 626
rect 665 625 666 626
rect 320 380 321 381
rect 322 380 323 381
rect 323 380 324 381
rect 325 380 326 381
rect 320 381 326 385
rect 320 385 321 386
rect 322 385 323 386
rect 323 385 324 386
rect 325 385 326 386
rect 580 800 581 801
rect 582 800 583 801
rect 583 800 584 801
rect 585 800 586 801
rect 580 801 586 805
rect 580 805 581 806
rect 582 805 583 806
rect 583 805 584 806
rect 585 805 586 806
rect 200 440 201 441
rect 202 440 203 441
rect 203 440 204 441
rect 205 440 206 441
rect 200 441 206 445
rect 200 445 201 446
rect 202 445 203 446
rect 203 445 204 446
rect 205 445 206 446
rect 320 580 321 581
rect 322 580 323 581
rect 323 580 324 581
rect 325 580 326 581
rect 320 581 326 585
rect 320 585 321 586
rect 322 585 323 586
rect 323 585 324 586
rect 325 585 326 586
rect 220 360 221 361
rect 222 360 223 361
rect 223 360 224 361
rect 225 360 226 361
rect 220 361 226 365
rect 220 365 221 366
rect 222 365 223 366
rect 223 365 224 366
rect 225 365 226 366
rect 260 340 261 341
rect 262 340 263 341
rect 263 340 264 341
rect 265 340 266 341
rect 260 341 266 345
rect 260 345 261 346
rect 262 345 263 346
rect 263 345 264 346
rect 265 345 266 346
rect 640 560 641 561
rect 642 560 643 561
rect 643 560 644 561
rect 645 560 646 561
rect 640 561 646 565
rect 640 565 641 566
rect 642 565 643 566
rect 643 565 644 566
rect 645 565 646 566
rect 160 440 161 441
rect 162 440 163 441
rect 163 440 164 441
rect 165 440 166 441
rect 160 441 166 445
rect 160 445 161 446
rect 162 445 163 446
rect 163 445 164 446
rect 165 445 166 446
rect 620 720 621 721
rect 622 720 623 721
rect 623 720 624 721
rect 625 720 626 721
rect 620 721 626 725
rect 620 725 621 726
rect 622 725 623 726
rect 623 725 624 726
rect 625 725 626 726
rect 460 720 461 721
rect 462 720 463 721
rect 463 720 464 721
rect 465 720 466 721
rect 460 721 466 725
rect 460 725 461 726
rect 462 725 463 726
rect 463 725 464 726
rect 465 725 466 726
rect 480 660 481 661
rect 482 660 483 661
rect 483 660 484 661
rect 485 660 486 661
rect 480 661 486 665
rect 480 665 481 666
rect 482 665 483 666
rect 483 665 484 666
rect 485 665 486 666
rect 600 460 601 461
rect 602 460 603 461
rect 603 460 604 461
rect 605 460 606 461
rect 600 461 606 465
rect 600 465 601 466
rect 602 465 603 466
rect 603 465 604 466
rect 605 465 606 466
rect 380 480 381 481
rect 382 480 383 481
rect 383 480 384 481
rect 385 480 386 481
rect 380 481 386 485
rect 380 485 381 486
rect 382 485 383 486
rect 383 485 384 486
rect 385 485 386 486
rect 720 680 721 681
rect 722 680 723 681
rect 723 680 724 681
rect 725 680 726 681
rect 720 681 726 685
rect 720 685 721 686
rect 722 685 723 686
rect 723 685 724 686
rect 725 685 726 686
rect 540 460 541 461
rect 542 460 543 461
rect 543 460 544 461
rect 545 460 546 461
rect 540 461 546 465
rect 540 465 541 466
rect 542 465 543 466
rect 543 465 544 466
rect 545 465 546 466
rect 620 500 621 501
rect 622 500 623 501
rect 623 500 624 501
rect 625 500 626 501
rect 620 501 626 505
rect 620 505 621 506
rect 622 505 623 506
rect 623 505 624 506
rect 625 505 626 506
rect 380 280 381 281
rect 382 280 383 281
rect 383 280 384 281
rect 385 280 386 281
rect 380 281 386 285
rect 380 285 381 286
rect 382 285 383 286
rect 383 285 384 286
rect 385 285 386 286
rect 820 660 821 661
rect 822 660 823 661
rect 823 660 824 661
rect 825 660 826 661
rect 820 661 826 665
rect 820 665 821 666
rect 822 665 823 666
rect 823 665 824 666
rect 825 665 826 666
rect 120 500 121 501
rect 122 500 123 501
rect 123 500 124 501
rect 125 500 126 501
rect 120 501 126 505
rect 120 505 121 506
rect 122 505 123 506
rect 123 505 124 506
rect 125 505 126 506
rect 500 800 501 801
rect 502 800 503 801
rect 503 800 504 801
rect 505 800 506 801
rect 500 801 506 805
rect 500 805 501 806
rect 502 805 503 806
rect 503 805 504 806
rect 505 805 506 806
rect 640 300 641 301
rect 642 300 643 301
rect 643 300 644 301
rect 645 300 646 301
rect 640 301 646 305
rect 640 305 641 306
rect 642 305 643 306
rect 643 305 644 306
rect 645 305 646 306
rect 800 460 801 461
rect 802 460 803 461
rect 803 460 804 461
rect 805 460 806 461
rect 800 461 806 465
rect 800 465 801 466
rect 802 465 803 466
rect 803 465 804 466
rect 805 465 806 466
rect 480 280 481 281
rect 482 280 483 281
rect 483 280 484 281
rect 485 280 486 281
rect 480 281 486 285
rect 480 285 481 286
rect 482 285 483 286
rect 483 285 484 286
rect 485 285 486 286
rect 740 700 741 701
rect 742 700 743 701
rect 743 700 744 701
rect 745 700 746 701
rect 740 701 746 705
rect 740 705 741 706
rect 742 705 743 706
rect 743 705 744 706
rect 745 705 746 706
rect 800 380 801 381
rect 802 380 803 381
rect 803 380 804 381
rect 805 380 806 381
rect 800 381 806 385
rect 800 385 801 386
rect 802 385 803 386
rect 803 385 804 386
rect 805 385 806 386
rect 420 680 421 681
rect 422 680 423 681
rect 423 680 424 681
rect 425 680 426 681
rect 420 681 426 685
rect 420 685 421 686
rect 422 685 423 686
rect 423 685 424 686
rect 425 685 426 686
rect 440 180 441 181
rect 442 180 443 181
rect 443 180 444 181
rect 445 180 446 181
rect 440 181 446 185
rect 440 185 441 186
rect 442 185 443 186
rect 443 185 444 186
rect 445 185 446 186
rect 500 840 501 841
rect 502 840 503 841
rect 503 840 504 841
rect 505 840 506 841
rect 500 841 506 845
rect 500 845 501 846
rect 502 845 503 846
rect 503 845 504 846
rect 505 845 506 846
rect 540 640 541 641
rect 542 640 543 641
rect 543 640 544 641
rect 545 640 546 641
rect 540 641 546 645
rect 540 645 541 646
rect 542 645 543 646
rect 543 645 544 646
rect 545 645 546 646
rect 620 260 621 261
rect 622 260 623 261
rect 623 260 624 261
rect 625 260 626 261
rect 620 261 626 265
rect 620 265 621 266
rect 622 265 623 266
rect 623 265 624 266
rect 625 265 626 266
rect 480 860 481 861
rect 482 860 483 861
rect 483 860 484 861
rect 485 860 486 861
rect 480 861 486 865
rect 480 865 481 866
rect 482 865 483 866
rect 483 865 484 866
rect 485 865 486 866
rect 440 800 441 801
rect 442 800 443 801
rect 443 800 444 801
rect 445 800 446 801
rect 440 801 446 805
rect 440 805 441 806
rect 442 805 443 806
rect 443 805 444 806
rect 445 805 446 806
rect 820 460 821 461
rect 822 460 823 461
rect 823 460 824 461
rect 825 460 826 461
rect 820 461 826 465
rect 820 465 821 466
rect 822 465 823 466
rect 823 465 824 466
rect 825 465 826 466
rect 600 740 601 741
rect 602 740 603 741
rect 603 740 604 741
rect 605 740 606 741
rect 600 741 606 745
rect 600 745 601 746
rect 602 745 603 746
rect 603 745 604 746
rect 605 745 606 746
rect 460 680 461 681
rect 462 680 463 681
rect 463 680 464 681
rect 465 680 466 681
rect 460 681 466 685
rect 460 685 461 686
rect 462 685 463 686
rect 463 685 464 686
rect 465 685 466 686
rect 220 480 221 481
rect 222 480 223 481
rect 223 480 224 481
rect 225 480 226 481
rect 220 481 226 485
rect 220 485 221 486
rect 222 485 223 486
rect 223 485 224 486
rect 225 485 226 486
rect 660 540 661 541
rect 662 540 663 541
rect 663 540 664 541
rect 665 540 666 541
rect 660 541 666 545
rect 660 545 661 546
rect 662 545 663 546
rect 663 545 664 546
rect 665 545 666 546
rect 340 720 341 721
rect 342 720 343 721
rect 343 720 344 721
rect 345 720 346 721
rect 340 721 346 725
rect 340 725 341 726
rect 342 725 343 726
rect 343 725 344 726
rect 345 725 346 726
rect 440 880 441 881
rect 442 880 443 881
rect 443 880 444 881
rect 445 880 446 881
rect 440 881 446 885
rect 440 885 441 886
rect 442 885 443 886
rect 443 885 444 886
rect 445 885 446 886
rect 400 800 401 801
rect 402 800 403 801
rect 403 800 404 801
rect 405 800 406 801
rect 400 801 406 805
rect 400 805 401 806
rect 402 805 403 806
rect 403 805 404 806
rect 405 805 406 806
rect 140 580 141 581
rect 142 580 143 581
rect 143 580 144 581
rect 145 580 146 581
rect 140 581 146 585
rect 140 585 141 586
rect 142 585 143 586
rect 143 585 144 586
rect 145 585 146 586
rect 180 580 181 581
rect 182 580 183 581
rect 183 580 184 581
rect 185 580 186 581
rect 180 581 186 585
rect 180 585 181 586
rect 182 585 183 586
rect 183 585 184 586
rect 185 585 186 586
rect 720 720 721 721
rect 722 720 723 721
rect 723 720 724 721
rect 725 720 726 721
rect 720 721 726 725
rect 720 725 721 726
rect 722 725 723 726
rect 723 725 724 726
rect 725 725 726 726
rect 320 480 321 481
rect 322 480 323 481
rect 323 480 324 481
rect 325 480 326 481
rect 320 481 326 485
rect 320 485 321 486
rect 322 485 323 486
rect 323 485 324 486
rect 325 485 326 486
rect 620 620 621 621
rect 622 620 623 621
rect 623 620 624 621
rect 625 620 626 621
rect 620 621 626 625
rect 620 625 621 626
rect 622 625 623 626
rect 623 625 624 626
rect 625 625 626 626
rect 560 800 561 801
rect 562 800 563 801
rect 563 800 564 801
rect 565 800 566 801
rect 560 801 566 805
rect 560 805 561 806
rect 562 805 563 806
rect 563 805 564 806
rect 565 805 566 806
rect 280 760 281 761
rect 282 760 283 761
rect 283 760 284 761
rect 285 760 286 761
rect 280 761 286 765
rect 280 765 281 766
rect 282 765 283 766
rect 283 765 284 766
rect 285 765 286 766
rect 800 680 801 681
rect 802 680 803 681
rect 803 680 804 681
rect 805 680 806 681
rect 800 681 806 685
rect 800 685 801 686
rect 802 685 803 686
rect 803 685 804 686
rect 805 685 806 686
rect 540 560 541 561
rect 542 560 543 561
rect 543 560 544 561
rect 545 560 546 561
rect 540 561 546 565
rect 540 565 541 566
rect 542 565 543 566
rect 543 565 544 566
rect 545 565 546 566
rect 440 500 441 501
rect 442 500 443 501
rect 443 500 444 501
rect 445 500 446 501
rect 440 501 446 505
rect 440 505 441 506
rect 442 505 443 506
rect 443 505 444 506
rect 445 505 446 506
rect 780 380 781 381
rect 782 380 783 381
rect 783 380 784 381
rect 785 380 786 381
rect 780 381 786 385
rect 780 385 781 386
rect 782 385 783 386
rect 783 385 784 386
rect 785 385 786 386
rect 800 600 801 601
rect 802 600 803 601
rect 803 600 804 601
rect 805 600 806 601
rect 800 601 806 605
rect 800 605 801 606
rect 802 605 803 606
rect 803 605 804 606
rect 805 605 806 606
rect 640 700 641 701
rect 642 700 643 701
rect 643 700 644 701
rect 645 700 646 701
rect 640 701 646 705
rect 640 705 641 706
rect 642 705 643 706
rect 643 705 644 706
rect 645 705 646 706
rect 500 760 501 761
rect 502 760 503 761
rect 503 760 504 761
rect 505 760 506 761
rect 500 761 506 765
rect 500 765 501 766
rect 502 765 503 766
rect 503 765 504 766
rect 505 765 506 766
rect 320 360 321 361
rect 322 360 323 361
rect 323 360 324 361
rect 325 360 326 361
rect 320 361 326 365
rect 320 365 321 366
rect 322 365 323 366
rect 323 365 324 366
rect 325 365 326 366
rect 160 560 161 561
rect 162 560 163 561
rect 163 560 164 561
rect 165 560 166 561
rect 160 561 166 565
rect 160 565 161 566
rect 162 565 163 566
rect 163 565 164 566
rect 165 565 166 566
rect 420 380 421 381
rect 422 380 423 381
rect 423 380 424 381
rect 425 380 426 381
rect 420 381 426 385
rect 420 385 421 386
rect 422 385 423 386
rect 423 385 424 386
rect 425 385 426 386
rect 140 620 141 621
rect 142 620 143 621
rect 143 620 144 621
rect 145 620 146 621
rect 140 621 146 625
rect 140 625 141 626
rect 142 625 143 626
rect 143 625 144 626
rect 145 625 146 626
rect 680 580 681 581
rect 682 580 683 581
rect 683 580 684 581
rect 685 580 686 581
rect 680 581 686 585
rect 680 585 681 586
rect 682 585 683 586
rect 683 585 684 586
rect 685 585 686 586
rect 780 620 781 621
rect 782 620 783 621
rect 783 620 784 621
rect 785 620 786 621
rect 780 621 786 625
rect 780 625 781 626
rect 782 625 783 626
rect 783 625 784 626
rect 785 625 786 626
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect 320 620 321 621
rect 322 620 323 621
rect 323 620 324 621
rect 325 620 326 621
rect 320 621 326 625
rect 320 625 321 626
rect 322 625 323 626
rect 323 625 324 626
rect 325 625 326 626
rect 720 440 721 441
rect 722 440 723 441
rect 723 440 724 441
rect 725 440 726 441
rect 720 441 726 445
rect 720 445 721 446
rect 722 445 723 446
rect 723 445 724 446
rect 725 445 726 446
rect 480 580 481 581
rect 482 580 483 581
rect 483 580 484 581
rect 485 580 486 581
rect 480 581 486 585
rect 480 585 481 586
rect 482 585 483 586
rect 483 585 484 586
rect 485 585 486 586
rect 340 740 341 741
rect 342 740 343 741
rect 343 740 344 741
rect 345 740 346 741
rect 340 741 346 745
rect 340 745 341 746
rect 342 745 343 746
rect 343 745 344 746
rect 345 745 346 746
rect 180 640 181 641
rect 182 640 183 641
rect 183 640 184 641
rect 185 640 186 641
rect 180 641 186 645
rect 180 645 181 646
rect 182 645 183 646
rect 183 645 184 646
rect 185 645 186 646
rect 800 440 801 441
rect 802 440 803 441
rect 803 440 804 441
rect 805 440 806 441
rect 800 441 806 445
rect 800 445 801 446
rect 802 445 803 446
rect 803 445 804 446
rect 805 445 806 446
rect 660 320 661 321
rect 662 320 663 321
rect 663 320 664 321
rect 665 320 666 321
rect 660 321 666 325
rect 660 325 661 326
rect 662 325 663 326
rect 663 325 664 326
rect 665 325 666 326
rect 260 740 261 741
rect 262 740 263 741
rect 263 740 264 741
rect 265 740 266 741
rect 260 741 266 745
rect 260 745 261 746
rect 262 745 263 746
rect 263 745 264 746
rect 265 745 266 746
rect 380 200 381 201
rect 382 200 383 201
rect 383 200 384 201
rect 385 200 386 201
rect 380 201 386 205
rect 380 205 381 206
rect 382 205 383 206
rect 383 205 384 206
rect 385 205 386 206
rect 620 380 621 381
rect 622 380 623 381
rect 623 380 624 381
rect 625 380 626 381
rect 620 381 626 385
rect 620 385 621 386
rect 622 385 623 386
rect 623 385 624 386
rect 625 385 626 386
rect 640 800 641 801
rect 642 800 643 801
rect 643 800 644 801
rect 645 800 646 801
rect 640 801 646 805
rect 640 805 641 806
rect 642 805 643 806
rect 643 805 644 806
rect 645 805 646 806
rect 480 160 481 161
rect 482 160 483 161
rect 483 160 484 161
rect 485 160 486 161
rect 480 161 486 165
rect 480 165 481 166
rect 482 165 483 166
rect 483 165 484 166
rect 485 165 486 166
rect 260 720 261 721
rect 262 720 263 721
rect 263 720 264 721
rect 265 720 266 721
rect 260 721 266 725
rect 260 725 261 726
rect 262 725 263 726
rect 263 725 264 726
rect 265 725 266 726
rect 580 480 581 481
rect 582 480 583 481
rect 583 480 584 481
rect 585 480 586 481
rect 580 481 586 485
rect 580 485 581 486
rect 582 485 583 486
rect 583 485 584 486
rect 585 485 586 486
rect 440 780 441 781
rect 442 780 443 781
rect 443 780 444 781
rect 445 780 446 781
rect 440 781 446 785
rect 440 785 441 786
rect 442 785 443 786
rect 443 785 444 786
rect 445 785 446 786
rect 860 500 861 501
rect 862 500 863 501
rect 863 500 864 501
rect 865 500 866 501
rect 860 501 866 505
rect 860 505 861 506
rect 862 505 863 506
rect 863 505 864 506
rect 865 505 866 506
rect 840 400 841 401
rect 842 400 843 401
rect 843 400 844 401
rect 845 400 846 401
rect 840 401 846 405
rect 840 405 841 406
rect 842 405 843 406
rect 843 405 844 406
rect 845 405 846 406
rect 320 600 321 601
rect 322 600 323 601
rect 323 600 324 601
rect 325 600 326 601
rect 320 601 326 605
rect 320 605 321 606
rect 322 605 323 606
rect 323 605 324 606
rect 325 605 326 606
rect 520 820 521 821
rect 522 820 523 821
rect 523 820 524 821
rect 525 820 526 821
rect 520 821 526 825
rect 520 825 521 826
rect 522 825 523 826
rect 523 825 524 826
rect 525 825 526 826
rect 520 860 521 861
rect 522 860 523 861
rect 523 860 524 861
rect 525 860 526 861
rect 520 861 526 865
rect 520 865 521 866
rect 522 865 523 866
rect 523 865 524 866
rect 525 865 526 866
rect 480 640 481 641
rect 482 640 483 641
rect 483 640 484 641
rect 485 640 486 641
rect 480 641 486 645
rect 480 645 481 646
rect 482 645 483 646
rect 483 645 484 646
rect 485 645 486 646
rect 720 500 721 501
rect 722 500 723 501
rect 723 500 724 501
rect 725 500 726 501
rect 720 501 726 505
rect 720 505 721 506
rect 722 505 723 506
rect 723 505 724 506
rect 725 505 726 506
rect 660 200 661 201
rect 662 200 663 201
rect 663 200 664 201
rect 665 200 666 201
rect 660 201 666 205
rect 660 205 661 206
rect 662 205 663 206
rect 663 205 664 206
rect 665 205 666 206
rect 400 420 401 421
rect 402 420 403 421
rect 403 420 404 421
rect 405 420 406 421
rect 400 421 406 425
rect 400 425 401 426
rect 402 425 403 426
rect 403 425 404 426
rect 405 425 406 426
rect 400 820 401 821
rect 402 820 403 821
rect 403 820 404 821
rect 405 820 406 821
rect 400 821 406 825
rect 400 825 401 826
rect 402 825 403 826
rect 403 825 404 826
rect 405 825 406 826
rect 740 300 741 301
rect 742 300 743 301
rect 743 300 744 301
rect 745 300 746 301
rect 740 301 746 305
rect 740 305 741 306
rect 742 305 743 306
rect 743 305 744 306
rect 745 305 746 306
rect 460 620 461 621
rect 462 620 463 621
rect 463 620 464 621
rect 465 620 466 621
rect 460 621 466 625
rect 460 625 461 626
rect 462 625 463 626
rect 463 625 464 626
rect 465 625 466 626
rect 620 700 621 701
rect 622 700 623 701
rect 623 700 624 701
rect 625 700 626 701
rect 620 701 626 705
rect 620 705 621 706
rect 622 705 623 706
rect 623 705 624 706
rect 625 705 626 706
rect 160 580 161 581
rect 162 580 163 581
rect 163 580 164 581
rect 165 580 166 581
rect 160 581 166 585
rect 160 585 161 586
rect 162 585 163 586
rect 163 585 164 586
rect 165 585 166 586
rect 460 660 461 661
rect 462 660 463 661
rect 463 660 464 661
rect 465 660 466 661
rect 460 661 466 665
rect 460 665 461 666
rect 462 665 463 666
rect 463 665 464 666
rect 465 665 466 666
rect 260 380 261 381
rect 262 380 263 381
rect 263 380 264 381
rect 265 380 266 381
rect 260 381 266 385
rect 260 385 261 386
rect 262 385 263 386
rect 263 385 264 386
rect 265 385 266 386
rect 560 640 561 641
rect 562 640 563 641
rect 563 640 564 641
rect 565 640 566 641
rect 560 641 566 645
rect 560 645 561 646
rect 562 645 563 646
rect 563 645 564 646
rect 565 645 566 646
rect 340 440 341 441
rect 342 440 343 441
rect 343 440 344 441
rect 345 440 346 441
rect 340 441 346 445
rect 340 445 341 446
rect 342 445 343 446
rect 343 445 344 446
rect 345 445 346 446
rect 280 300 281 301
rect 282 300 283 301
rect 283 300 284 301
rect 285 300 286 301
rect 280 301 286 305
rect 280 305 281 306
rect 282 305 283 306
rect 283 305 284 306
rect 285 305 286 306
rect 400 260 401 261
rect 402 260 403 261
rect 403 260 404 261
rect 405 260 406 261
rect 400 261 406 265
rect 400 265 401 266
rect 402 265 403 266
rect 403 265 404 266
rect 405 265 406 266
rect 500 860 501 861
rect 502 860 503 861
rect 503 860 504 861
rect 505 860 506 861
rect 500 861 506 865
rect 500 865 501 866
rect 502 865 503 866
rect 503 865 504 866
rect 505 865 506 866
rect 400 220 401 221
rect 402 220 403 221
rect 403 220 404 221
rect 405 220 406 221
rect 400 221 406 225
rect 400 225 401 226
rect 402 225 403 226
rect 403 225 404 226
rect 405 225 406 226
rect 360 220 361 221
rect 362 220 363 221
rect 363 220 364 221
rect 365 220 366 221
rect 360 221 366 225
rect 360 225 361 226
rect 362 225 363 226
rect 363 225 364 226
rect 365 225 366 226
rect 760 480 761 481
rect 762 480 763 481
rect 763 480 764 481
rect 765 480 766 481
rect 760 481 766 485
rect 760 485 761 486
rect 762 485 763 486
rect 763 485 764 486
rect 765 485 766 486
rect 640 500 641 501
rect 642 500 643 501
rect 643 500 644 501
rect 645 500 646 501
rect 640 501 646 505
rect 640 505 641 506
rect 642 505 643 506
rect 643 505 644 506
rect 645 505 646 506
rect 520 580 521 581
rect 522 580 523 581
rect 523 580 524 581
rect 525 580 526 581
rect 520 581 526 585
rect 520 585 521 586
rect 522 585 523 586
rect 523 585 524 586
rect 525 585 526 586
rect 380 520 381 521
rect 382 520 383 521
rect 383 520 384 521
rect 385 520 386 521
rect 380 521 386 525
rect 380 525 381 526
rect 382 525 383 526
rect 383 525 384 526
rect 385 525 386 526
rect 460 440 461 441
rect 462 440 463 441
rect 463 440 464 441
rect 465 440 466 441
rect 460 441 466 445
rect 460 445 461 446
rect 462 445 463 446
rect 463 445 464 446
rect 465 445 466 446
rect 780 360 781 361
rect 782 360 783 361
rect 783 360 784 361
rect 785 360 786 361
rect 780 361 786 365
rect 780 365 781 366
rect 782 365 783 366
rect 783 365 784 366
rect 785 365 786 366
rect 540 900 541 901
rect 542 900 543 901
rect 543 900 544 901
rect 545 900 546 901
rect 540 901 546 905
rect 540 905 541 906
rect 542 905 543 906
rect 543 905 544 906
rect 545 905 546 906
rect 360 800 361 801
rect 362 800 363 801
rect 363 800 364 801
rect 365 800 366 801
rect 360 801 366 805
rect 360 805 361 806
rect 362 805 363 806
rect 363 805 364 806
rect 365 805 366 806
rect 180 540 181 541
rect 182 540 183 541
rect 183 540 184 541
rect 185 540 186 541
rect 180 541 186 545
rect 180 545 181 546
rect 182 545 183 546
rect 183 545 184 546
rect 185 545 186 546
rect 260 500 261 501
rect 262 500 263 501
rect 263 500 264 501
rect 265 500 266 501
rect 260 501 266 505
rect 260 505 261 506
rect 262 505 263 506
rect 263 505 264 506
rect 265 505 266 506
rect 380 720 381 721
rect 382 720 383 721
rect 383 720 384 721
rect 385 720 386 721
rect 380 721 386 725
rect 380 725 381 726
rect 382 725 383 726
rect 383 725 384 726
rect 385 725 386 726
rect 480 300 481 301
rect 482 300 483 301
rect 483 300 484 301
rect 485 300 486 301
rect 480 301 486 305
rect 480 305 481 306
rect 482 305 483 306
rect 483 305 484 306
rect 485 305 486 306
rect 300 380 301 381
rect 302 380 303 381
rect 303 380 304 381
rect 305 380 306 381
rect 300 381 306 385
rect 300 385 301 386
rect 302 385 303 386
rect 303 385 304 386
rect 305 385 306 386
rect 420 200 421 201
rect 422 200 423 201
rect 423 200 424 201
rect 425 200 426 201
rect 420 201 426 205
rect 420 205 421 206
rect 422 205 423 206
rect 423 205 424 206
rect 425 205 426 206
rect 580 200 581 201
rect 582 200 583 201
rect 583 200 584 201
rect 585 200 586 201
rect 580 201 586 205
rect 580 205 581 206
rect 582 205 583 206
rect 583 205 584 206
rect 585 205 586 206
rect 560 660 561 661
rect 562 660 563 661
rect 563 660 564 661
rect 565 660 566 661
rect 560 661 566 665
rect 560 665 561 666
rect 562 665 563 666
rect 563 665 564 666
rect 565 665 566 666
rect 640 840 641 841
rect 642 840 643 841
rect 643 840 644 841
rect 645 840 646 841
rect 640 841 646 845
rect 640 845 641 846
rect 642 845 643 846
rect 643 845 644 846
rect 645 845 646 846
rect 420 600 421 601
rect 422 600 423 601
rect 423 600 424 601
rect 425 600 426 601
rect 420 601 426 605
rect 420 605 421 606
rect 422 605 423 606
rect 423 605 424 606
rect 425 605 426 606
rect 280 500 281 501
rect 282 500 283 501
rect 283 500 284 501
rect 285 500 286 501
rect 280 501 286 505
rect 280 505 281 506
rect 282 505 283 506
rect 283 505 284 506
rect 285 505 286 506
rect 420 400 421 401
rect 422 400 423 401
rect 423 400 424 401
rect 425 400 426 401
rect 420 401 426 405
rect 420 405 421 406
rect 422 405 423 406
rect 423 405 424 406
rect 425 405 426 406
rect 680 400 681 401
rect 682 400 683 401
rect 683 400 684 401
rect 685 400 686 401
rect 680 401 686 405
rect 680 405 681 406
rect 682 405 683 406
rect 683 405 684 406
rect 685 405 686 406
rect 240 380 241 381
rect 242 380 243 381
rect 243 380 244 381
rect 245 380 246 381
rect 240 381 246 385
rect 240 385 241 386
rect 242 385 243 386
rect 243 385 244 386
rect 245 385 246 386
rect 320 640 321 641
rect 322 640 323 641
rect 323 640 324 641
rect 325 640 326 641
rect 320 641 326 645
rect 320 645 321 646
rect 322 645 323 646
rect 323 645 324 646
rect 325 645 326 646
rect 320 340 321 341
rect 322 340 323 341
rect 323 340 324 341
rect 325 340 326 341
rect 320 341 326 345
rect 320 345 321 346
rect 322 345 323 346
rect 323 345 324 346
rect 325 345 326 346
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect 400 540 401 541
rect 402 540 403 541
rect 403 540 404 541
rect 405 540 406 541
rect 400 541 406 545
rect 400 545 401 546
rect 402 545 403 546
rect 403 545 404 546
rect 405 545 406 546
rect 300 480 301 481
rect 302 480 303 481
rect 303 480 304 481
rect 305 480 306 481
rect 300 481 306 485
rect 300 485 301 486
rect 302 485 303 486
rect 303 485 304 486
rect 305 485 306 486
rect 420 340 421 341
rect 422 340 423 341
rect 423 340 424 341
rect 425 340 426 341
rect 420 341 426 345
rect 420 345 421 346
rect 422 345 423 346
rect 423 345 424 346
rect 425 345 426 346
rect 820 520 821 521
rect 822 520 823 521
rect 823 520 824 521
rect 825 520 826 521
rect 820 521 826 525
rect 820 525 821 526
rect 822 525 823 526
rect 823 525 824 526
rect 825 525 826 526
rect 200 660 201 661
rect 202 660 203 661
rect 203 660 204 661
rect 205 660 206 661
rect 200 661 206 665
rect 200 665 201 666
rect 202 665 203 666
rect 203 665 204 666
rect 205 665 206 666
rect 600 420 601 421
rect 602 420 603 421
rect 603 420 604 421
rect 605 420 606 421
rect 600 421 606 425
rect 600 425 601 426
rect 602 425 603 426
rect 603 425 604 426
rect 605 425 606 426
rect 820 580 821 581
rect 822 580 823 581
rect 823 580 824 581
rect 825 580 826 581
rect 820 581 826 585
rect 820 585 821 586
rect 822 585 823 586
rect 823 585 824 586
rect 825 585 826 586
rect 360 340 361 341
rect 362 340 363 341
rect 363 340 364 341
rect 365 340 366 341
rect 360 341 366 345
rect 360 345 361 346
rect 362 345 363 346
rect 363 345 364 346
rect 365 345 366 346
rect 640 540 641 541
rect 642 540 643 541
rect 643 540 644 541
rect 645 540 646 541
rect 640 541 646 545
rect 640 545 641 546
rect 642 545 643 546
rect 643 545 644 546
rect 645 545 646 546
rect 640 340 641 341
rect 642 340 643 341
rect 643 340 644 341
rect 645 340 646 341
rect 640 341 646 345
rect 640 345 641 346
rect 642 345 643 346
rect 643 345 644 346
rect 645 345 646 346
rect 480 460 481 461
rect 482 460 483 461
rect 483 460 484 461
rect 485 460 486 461
rect 480 461 486 465
rect 480 465 481 466
rect 482 465 483 466
rect 483 465 484 466
rect 485 465 486 466
rect 480 340 481 341
rect 482 340 483 341
rect 483 340 484 341
rect 485 340 486 341
rect 480 341 486 345
rect 480 345 481 346
rect 482 345 483 346
rect 483 345 484 346
rect 485 345 486 346
rect 360 440 361 441
rect 362 440 363 441
rect 363 440 364 441
rect 365 440 366 441
rect 360 441 366 445
rect 360 445 361 446
rect 362 445 363 446
rect 363 445 364 446
rect 365 445 366 446
rect 660 340 661 341
rect 662 340 663 341
rect 663 340 664 341
rect 665 340 666 341
rect 660 341 666 345
rect 660 345 661 346
rect 662 345 663 346
rect 663 345 664 346
rect 665 345 666 346
rect 280 740 281 741
rect 282 740 283 741
rect 283 740 284 741
rect 285 740 286 741
rect 280 741 286 745
rect 280 745 281 746
rect 282 745 283 746
rect 283 745 284 746
rect 285 745 286 746
rect 700 500 701 501
rect 702 500 703 501
rect 703 500 704 501
rect 705 500 706 501
rect 700 501 706 505
rect 700 505 701 506
rect 702 505 703 506
rect 703 505 704 506
rect 705 505 706 506
rect 260 320 261 321
rect 262 320 263 321
rect 263 320 264 321
rect 265 320 266 321
rect 260 321 266 325
rect 260 325 261 326
rect 262 325 263 326
rect 263 325 264 326
rect 265 325 266 326
rect 380 340 381 341
rect 382 340 383 341
rect 383 340 384 341
rect 385 340 386 341
rect 380 341 386 345
rect 380 345 381 346
rect 382 345 383 346
rect 383 345 384 346
rect 385 345 386 346
rect 700 540 701 541
rect 702 540 703 541
rect 703 540 704 541
rect 705 540 706 541
rect 700 541 706 545
rect 700 545 701 546
rect 702 545 703 546
rect 703 545 704 546
rect 705 545 706 546
rect 880 520 881 521
rect 882 520 883 521
rect 883 520 884 521
rect 885 520 886 521
rect 880 521 886 525
rect 880 525 881 526
rect 882 525 883 526
rect 883 525 884 526
rect 885 525 886 526
rect 840 540 841 541
rect 842 540 843 541
rect 843 540 844 541
rect 845 540 846 541
rect 840 541 846 545
rect 840 545 841 546
rect 842 545 843 546
rect 843 545 844 546
rect 845 545 846 546
rect 620 780 621 781
rect 622 780 623 781
rect 623 780 624 781
rect 625 780 626 781
rect 620 781 626 785
rect 620 785 621 786
rect 622 785 623 786
rect 623 785 624 786
rect 625 785 626 786
rect 320 540 321 541
rect 322 540 323 541
rect 323 540 324 541
rect 325 540 326 541
rect 320 541 326 545
rect 320 545 321 546
rect 322 545 323 546
rect 323 545 324 546
rect 325 545 326 546
rect 760 700 761 701
rect 762 700 763 701
rect 763 700 764 701
rect 765 700 766 701
rect 760 701 766 705
rect 760 705 761 706
rect 762 705 763 706
rect 763 705 764 706
rect 765 705 766 706
rect 360 780 361 781
rect 362 780 363 781
rect 363 780 364 781
rect 365 780 366 781
rect 360 781 366 785
rect 360 785 361 786
rect 362 785 363 786
rect 363 785 364 786
rect 365 785 366 786
rect 420 820 421 821
rect 422 820 423 821
rect 423 820 424 821
rect 425 820 426 821
rect 420 821 426 825
rect 420 825 421 826
rect 422 825 423 826
rect 423 825 424 826
rect 425 825 426 826
rect 740 720 741 721
rect 742 720 743 721
rect 743 720 744 721
rect 745 720 746 721
rect 740 721 746 725
rect 740 725 741 726
rect 742 725 743 726
rect 743 725 744 726
rect 745 725 746 726
rect 680 600 681 601
rect 682 600 683 601
rect 683 600 684 601
rect 685 600 686 601
rect 680 601 686 605
rect 680 605 681 606
rect 682 605 683 606
rect 683 605 684 606
rect 685 605 686 606
rect 640 220 641 221
rect 642 220 643 221
rect 643 220 644 221
rect 645 220 646 221
rect 640 221 646 225
rect 640 225 641 226
rect 642 225 643 226
rect 643 225 644 226
rect 645 225 646 226
rect 640 320 641 321
rect 642 320 643 321
rect 643 320 644 321
rect 645 320 646 321
rect 640 321 646 325
rect 640 325 641 326
rect 642 325 643 326
rect 643 325 644 326
rect 645 325 646 326
rect 780 640 781 641
rect 782 640 783 641
rect 783 640 784 641
rect 785 640 786 641
rect 780 641 786 645
rect 780 645 781 646
rect 782 645 783 646
rect 783 645 784 646
rect 785 645 786 646
rect 800 620 801 621
rect 802 620 803 621
rect 803 620 804 621
rect 805 620 806 621
rect 800 621 806 625
rect 800 625 801 626
rect 802 625 803 626
rect 803 625 804 626
rect 805 625 806 626
rect 460 220 461 221
rect 462 220 463 221
rect 463 220 464 221
rect 465 220 466 221
rect 460 221 466 225
rect 460 225 461 226
rect 462 225 463 226
rect 463 225 464 226
rect 465 225 466 226
rect 500 520 501 521
rect 502 520 503 521
rect 503 520 504 521
rect 505 520 506 521
rect 500 521 506 525
rect 500 525 501 526
rect 502 525 503 526
rect 503 525 504 526
rect 505 525 506 526
rect 440 300 441 301
rect 442 300 443 301
rect 443 300 444 301
rect 445 300 446 301
rect 440 301 446 305
rect 440 305 441 306
rect 442 305 443 306
rect 443 305 444 306
rect 445 305 446 306
rect 100 460 101 461
rect 102 460 103 461
rect 103 460 104 461
rect 105 460 106 461
rect 100 461 106 465
rect 100 465 101 466
rect 102 465 103 466
rect 103 465 104 466
rect 105 465 106 466
rect 180 520 181 521
rect 182 520 183 521
rect 183 520 184 521
rect 185 520 186 521
rect 180 521 186 525
rect 180 525 181 526
rect 182 525 183 526
rect 183 525 184 526
rect 185 525 186 526
rect 260 560 261 561
rect 262 560 263 561
rect 263 560 264 561
rect 265 560 266 561
rect 260 561 266 565
rect 260 565 261 566
rect 262 565 263 566
rect 263 565 264 566
rect 265 565 266 566
rect 600 400 601 401
rect 602 400 603 401
rect 603 400 604 401
rect 605 400 606 401
rect 600 401 606 405
rect 600 405 601 406
rect 602 405 603 406
rect 603 405 604 406
rect 605 405 606 406
rect 520 660 521 661
rect 522 660 523 661
rect 523 660 524 661
rect 525 660 526 661
rect 520 661 526 665
rect 520 665 521 666
rect 522 665 523 666
rect 523 665 524 666
rect 525 665 526 666
rect 140 520 141 521
rect 142 520 143 521
rect 143 520 144 521
rect 145 520 146 521
rect 140 521 146 525
rect 140 525 141 526
rect 142 525 143 526
rect 143 525 144 526
rect 145 525 146 526
rect 800 400 801 401
rect 802 400 803 401
rect 803 400 804 401
rect 805 400 806 401
rect 800 401 806 405
rect 800 405 801 406
rect 802 405 803 406
rect 803 405 804 406
rect 805 405 806 406
rect 580 820 581 821
rect 582 820 583 821
rect 583 820 584 821
rect 585 820 586 821
rect 580 821 586 825
rect 580 825 581 826
rect 582 825 583 826
rect 583 825 584 826
rect 585 825 586 826
rect 560 540 561 541
rect 562 540 563 541
rect 563 540 564 541
rect 565 540 566 541
rect 560 541 566 545
rect 560 545 561 546
rect 562 545 563 546
rect 563 545 564 546
rect 565 545 566 546
rect 200 500 201 501
rect 202 500 203 501
rect 203 500 204 501
rect 205 500 206 501
rect 200 501 206 505
rect 200 505 201 506
rect 202 505 203 506
rect 203 505 204 506
rect 205 505 206 506
rect 700 340 701 341
rect 702 340 703 341
rect 703 340 704 341
rect 705 340 706 341
rect 700 341 706 345
rect 700 345 701 346
rect 702 345 703 346
rect 703 345 704 346
rect 705 345 706 346
rect 560 420 561 421
rect 562 420 563 421
rect 563 420 564 421
rect 565 420 566 421
rect 560 421 566 425
rect 560 425 561 426
rect 562 425 563 426
rect 563 425 564 426
rect 565 425 566 426
rect 140 600 141 601
rect 142 600 143 601
rect 143 600 144 601
rect 145 600 146 601
rect 140 601 146 605
rect 140 605 141 606
rect 142 605 143 606
rect 143 605 144 606
rect 145 605 146 606
rect 500 380 501 381
rect 502 380 503 381
rect 503 380 504 381
rect 505 380 506 381
rect 500 381 506 385
rect 500 385 501 386
rect 502 385 503 386
rect 503 385 504 386
rect 505 385 506 386
rect 600 800 601 801
rect 602 800 603 801
rect 603 800 604 801
rect 605 800 606 801
rect 600 801 606 805
rect 600 805 601 806
rect 602 805 603 806
rect 603 805 604 806
rect 605 805 606 806
rect 440 620 441 621
rect 442 620 443 621
rect 443 620 444 621
rect 445 620 446 621
rect 440 621 446 625
rect 440 625 441 626
rect 442 625 443 626
rect 443 625 444 626
rect 445 625 446 626
rect 200 540 201 541
rect 202 540 203 541
rect 203 540 204 541
rect 205 540 206 541
rect 200 541 206 545
rect 200 545 201 546
rect 202 545 203 546
rect 203 545 204 546
rect 205 545 206 546
rect 160 420 161 421
rect 162 420 163 421
rect 163 420 164 421
rect 165 420 166 421
rect 160 421 166 425
rect 160 425 161 426
rect 162 425 163 426
rect 163 425 164 426
rect 165 425 166 426
rect 560 160 561 161
rect 562 160 563 161
rect 563 160 564 161
rect 565 160 566 161
rect 560 161 566 165
rect 560 165 561 166
rect 562 165 563 166
rect 563 165 564 166
rect 565 165 566 166
rect 380 760 381 761
rect 382 760 383 761
rect 383 760 384 761
rect 385 760 386 761
rect 380 761 386 765
rect 380 765 381 766
rect 382 765 383 766
rect 383 765 384 766
rect 385 765 386 766
rect 900 560 901 561
rect 902 560 903 561
rect 903 560 904 561
rect 905 560 906 561
rect 900 561 906 565
rect 900 565 901 566
rect 902 565 903 566
rect 903 565 904 566
rect 905 565 906 566
rect 280 600 281 601
rect 282 600 283 601
rect 283 600 284 601
rect 285 600 286 601
rect 280 601 286 605
rect 280 605 281 606
rect 282 605 283 606
rect 283 605 284 606
rect 285 605 286 606
rect 520 520 521 521
rect 522 520 523 521
rect 523 520 524 521
rect 525 520 526 521
rect 520 521 526 525
rect 520 525 521 526
rect 522 525 523 526
rect 523 525 524 526
rect 525 525 526 526
rect 520 420 521 421
rect 522 420 523 421
rect 523 420 524 421
rect 525 420 526 421
rect 520 421 526 425
rect 520 425 521 426
rect 522 425 523 426
rect 523 425 524 426
rect 525 425 526 426
rect 340 260 341 261
rect 342 260 343 261
rect 343 260 344 261
rect 345 260 346 261
rect 340 261 346 265
rect 340 265 341 266
rect 342 265 343 266
rect 343 265 344 266
rect 345 265 346 266
rect 200 520 201 521
rect 202 520 203 521
rect 203 520 204 521
rect 205 520 206 521
rect 200 521 206 525
rect 200 525 201 526
rect 202 525 203 526
rect 203 525 204 526
rect 205 525 206 526
rect 760 500 761 501
rect 762 500 763 501
rect 763 500 764 501
rect 765 500 766 501
rect 760 501 766 505
rect 760 505 761 506
rect 762 505 763 506
rect 763 505 764 506
rect 765 505 766 506
rect 880 500 881 501
rect 882 500 883 501
rect 883 500 884 501
rect 885 500 886 501
rect 880 501 886 505
rect 880 505 881 506
rect 882 505 883 506
rect 883 505 884 506
rect 885 505 886 506
rect 360 760 361 761
rect 362 760 363 761
rect 363 760 364 761
rect 365 760 366 761
rect 360 761 366 765
rect 360 765 361 766
rect 362 765 363 766
rect 363 765 364 766
rect 365 765 366 766
rect 580 780 581 781
rect 582 780 583 781
rect 583 780 584 781
rect 585 780 586 781
rect 580 781 586 785
rect 580 785 581 786
rect 582 785 583 786
rect 583 785 584 786
rect 585 785 586 786
rect 620 180 621 181
rect 622 180 623 181
rect 623 180 624 181
rect 625 180 626 181
rect 620 181 626 185
rect 620 185 621 186
rect 622 185 623 186
rect 623 185 624 186
rect 625 185 626 186
rect 340 400 341 401
rect 342 400 343 401
rect 343 400 344 401
rect 345 400 346 401
rect 340 401 346 405
rect 340 405 341 406
rect 342 405 343 406
rect 343 405 344 406
rect 345 405 346 406
rect 440 540 441 541
rect 442 540 443 541
rect 443 540 444 541
rect 445 540 446 541
rect 440 541 446 545
rect 440 545 441 546
rect 442 545 443 546
rect 443 545 444 546
rect 445 545 446 546
rect 820 600 821 601
rect 822 600 823 601
rect 823 600 824 601
rect 825 600 826 601
rect 820 601 826 605
rect 820 605 821 606
rect 822 605 823 606
rect 823 605 824 606
rect 825 605 826 606
rect 360 280 361 281
rect 362 280 363 281
rect 363 280 364 281
rect 365 280 366 281
rect 360 281 366 285
rect 360 285 361 286
rect 362 285 363 286
rect 363 285 364 286
rect 365 285 366 286
rect 540 500 541 501
rect 542 500 543 501
rect 543 500 544 501
rect 545 500 546 501
rect 540 501 546 505
rect 540 505 541 506
rect 542 505 543 506
rect 543 505 544 506
rect 545 505 546 506
rect 540 180 541 181
rect 542 180 543 181
rect 543 180 544 181
rect 545 180 546 181
rect 540 181 546 185
rect 540 185 541 186
rect 542 185 543 186
rect 543 185 544 186
rect 545 185 546 186
rect 400 760 401 761
rect 402 760 403 761
rect 403 760 404 761
rect 405 760 406 761
rect 400 761 406 765
rect 400 765 401 766
rect 402 765 403 766
rect 403 765 404 766
rect 405 765 406 766
rect 700 300 701 301
rect 702 300 703 301
rect 703 300 704 301
rect 705 300 706 301
rect 700 301 706 305
rect 700 305 701 306
rect 702 305 703 306
rect 703 305 704 306
rect 705 305 706 306
rect 280 540 281 541
rect 282 540 283 541
rect 283 540 284 541
rect 285 540 286 541
rect 280 541 286 545
rect 280 545 281 546
rect 282 545 283 546
rect 283 545 284 546
rect 285 545 286 546
rect 780 680 781 681
rect 782 680 783 681
rect 783 680 784 681
rect 785 680 786 681
rect 780 681 786 685
rect 780 685 781 686
rect 782 685 783 686
rect 783 685 784 686
rect 785 685 786 686
rect 180 660 181 661
rect 182 660 183 661
rect 183 660 184 661
rect 185 660 186 661
rect 180 661 186 665
rect 180 665 181 666
rect 182 665 183 666
rect 183 665 184 666
rect 185 665 186 666
rect 440 240 441 241
rect 442 240 443 241
rect 443 240 444 241
rect 445 240 446 241
rect 440 241 446 245
rect 440 245 441 246
rect 442 245 443 246
rect 443 245 444 246
rect 445 245 446 246
rect 340 820 341 821
rect 342 820 343 821
rect 343 820 344 821
rect 345 820 346 821
rect 340 821 346 825
rect 340 825 341 826
rect 342 825 343 826
rect 343 825 344 826
rect 345 825 346 826
rect 580 320 581 321
rect 582 320 583 321
rect 583 320 584 321
rect 585 320 586 321
rect 580 321 586 325
rect 580 325 581 326
rect 582 325 583 326
rect 583 325 584 326
rect 585 325 586 326
rect 320 720 321 721
rect 322 720 323 721
rect 323 720 324 721
rect 325 720 326 721
rect 320 721 326 725
rect 320 725 321 726
rect 322 725 323 726
rect 323 725 324 726
rect 325 725 326 726
rect 500 580 501 581
rect 502 580 503 581
rect 503 580 504 581
rect 505 580 506 581
rect 500 581 506 585
rect 500 585 501 586
rect 502 585 503 586
rect 503 585 504 586
rect 505 585 506 586
rect 540 140 541 141
rect 542 140 543 141
rect 543 140 544 141
rect 545 140 546 141
rect 540 141 546 145
rect 540 145 541 146
rect 542 145 543 146
rect 543 145 544 146
rect 545 145 546 146
rect 400 560 401 561
rect 402 560 403 561
rect 403 560 404 561
rect 405 560 406 561
rect 400 561 406 565
rect 400 565 401 566
rect 402 565 403 566
rect 403 565 404 566
rect 405 565 406 566
rect 660 500 661 501
rect 662 500 663 501
rect 663 500 664 501
rect 665 500 666 501
rect 660 501 666 505
rect 660 505 661 506
rect 662 505 663 506
rect 663 505 664 506
rect 665 505 666 506
rect 200 620 201 621
rect 202 620 203 621
rect 203 620 204 621
rect 205 620 206 621
rect 200 621 206 625
rect 200 625 201 626
rect 202 625 203 626
rect 203 625 204 626
rect 205 625 206 626
rect 580 760 581 761
rect 582 760 583 761
rect 583 760 584 761
rect 585 760 586 761
rect 580 761 586 765
rect 580 765 581 766
rect 582 765 583 766
rect 583 765 584 766
rect 585 765 586 766
rect 120 440 121 441
rect 122 440 123 441
rect 123 440 124 441
rect 125 440 126 441
rect 120 441 126 445
rect 120 445 121 446
rect 122 445 123 446
rect 123 445 124 446
rect 125 445 126 446
rect 480 840 481 841
rect 482 840 483 841
rect 483 840 484 841
rect 485 840 486 841
rect 480 841 486 845
rect 480 845 481 846
rect 482 845 483 846
rect 483 845 484 846
rect 485 845 486 846
rect 480 760 481 761
rect 482 760 483 761
rect 483 760 484 761
rect 485 760 486 761
rect 480 761 486 765
rect 480 765 481 766
rect 482 765 483 766
rect 483 765 484 766
rect 485 765 486 766
rect 300 420 301 421
rect 302 420 303 421
rect 303 420 304 421
rect 305 420 306 421
rect 300 421 306 425
rect 300 425 301 426
rect 302 425 303 426
rect 303 425 304 426
rect 305 425 306 426
rect 820 640 821 641
rect 822 640 823 641
rect 823 640 824 641
rect 825 640 826 641
rect 820 641 826 645
rect 820 645 821 646
rect 822 645 823 646
rect 823 645 824 646
rect 825 645 826 646
rect 520 560 521 561
rect 522 560 523 561
rect 523 560 524 561
rect 525 560 526 561
rect 520 561 526 565
rect 520 565 521 566
rect 522 565 523 566
rect 523 565 524 566
rect 525 565 526 566
rect 500 880 501 881
rect 502 880 503 881
rect 503 880 504 881
rect 505 880 506 881
rect 500 881 506 885
rect 500 885 501 886
rect 502 885 503 886
rect 503 885 504 886
rect 505 885 506 886
rect 320 500 321 501
rect 322 500 323 501
rect 323 500 324 501
rect 325 500 326 501
rect 320 501 326 505
rect 320 505 321 506
rect 322 505 323 506
rect 323 505 324 506
rect 325 505 326 506
rect 880 460 881 461
rect 882 460 883 461
rect 883 460 884 461
rect 885 460 886 461
rect 880 461 886 465
rect 880 465 881 466
rect 882 465 883 466
rect 883 465 884 466
rect 885 465 886 466
rect 580 220 581 221
rect 582 220 583 221
rect 583 220 584 221
rect 585 220 586 221
rect 580 221 586 225
rect 580 225 581 226
rect 582 225 583 226
rect 583 225 584 226
rect 585 225 586 226
rect 800 640 801 641
rect 802 640 803 641
rect 803 640 804 641
rect 805 640 806 641
rect 800 641 806 645
rect 800 645 801 646
rect 802 645 803 646
rect 803 645 804 646
rect 805 645 806 646
rect 160 520 161 521
rect 162 520 163 521
rect 163 520 164 521
rect 165 520 166 521
rect 160 521 166 525
rect 160 525 161 526
rect 162 525 163 526
rect 163 525 164 526
rect 165 525 166 526
rect 640 580 641 581
rect 642 580 643 581
rect 643 580 644 581
rect 645 580 646 581
rect 640 581 646 585
rect 640 585 641 586
rect 642 585 643 586
rect 643 585 644 586
rect 645 585 646 586
rect 540 320 541 321
rect 542 320 543 321
rect 543 320 544 321
rect 545 320 546 321
rect 540 321 546 325
rect 540 325 541 326
rect 542 325 543 326
rect 543 325 544 326
rect 545 325 546 326
rect 280 440 281 441
rect 282 440 283 441
rect 283 440 284 441
rect 285 440 286 441
rect 280 441 286 445
rect 280 445 281 446
rect 282 445 283 446
rect 283 445 284 446
rect 285 445 286 446
rect 600 840 601 841
rect 602 840 603 841
rect 603 840 604 841
rect 605 840 606 841
rect 600 841 606 845
rect 600 845 601 846
rect 602 845 603 846
rect 603 845 604 846
rect 605 845 606 846
rect 800 500 801 501
rect 802 500 803 501
rect 803 500 804 501
rect 805 500 806 501
rect 800 501 806 505
rect 800 505 801 506
rect 802 505 803 506
rect 803 505 804 506
rect 805 505 806 506
rect 300 720 301 721
rect 302 720 303 721
rect 303 720 304 721
rect 305 720 306 721
rect 300 721 306 725
rect 300 725 301 726
rect 302 725 303 726
rect 303 725 304 726
rect 305 725 306 726
rect 680 520 681 521
rect 682 520 683 521
rect 683 520 684 521
rect 685 520 686 521
rect 680 521 686 525
rect 680 525 681 526
rect 682 525 683 526
rect 683 525 684 526
rect 685 525 686 526
rect 420 840 421 841
rect 422 840 423 841
rect 423 840 424 841
rect 425 840 426 841
rect 420 841 426 845
rect 420 845 421 846
rect 422 845 423 846
rect 423 845 424 846
rect 425 845 426 846
rect 400 440 401 441
rect 402 440 403 441
rect 403 440 404 441
rect 405 440 406 441
rect 400 441 406 445
rect 400 445 401 446
rect 402 445 403 446
rect 403 445 404 446
rect 405 445 406 446
rect 440 360 441 361
rect 442 360 443 361
rect 443 360 444 361
rect 445 360 446 361
rect 440 361 446 365
rect 440 365 441 366
rect 442 365 443 366
rect 443 365 444 366
rect 445 365 446 366
rect 840 460 841 461
rect 842 460 843 461
rect 843 460 844 461
rect 845 460 846 461
rect 840 461 846 465
rect 840 465 841 466
rect 842 465 843 466
rect 843 465 844 466
rect 845 465 846 466
rect 300 740 301 741
rect 302 740 303 741
rect 303 740 304 741
rect 305 740 306 741
rect 300 741 306 745
rect 300 745 301 746
rect 302 745 303 746
rect 303 745 304 746
rect 305 745 306 746
rect 280 720 281 721
rect 282 720 283 721
rect 283 720 284 721
rect 285 720 286 721
rect 280 721 286 725
rect 280 725 281 726
rect 282 725 283 726
rect 283 725 284 726
rect 285 725 286 726
rect 380 600 381 601
rect 382 600 383 601
rect 383 600 384 601
rect 385 600 386 601
rect 380 601 386 605
rect 380 605 381 606
rect 382 605 383 606
rect 383 605 384 606
rect 385 605 386 606
rect 600 820 601 821
rect 602 820 603 821
rect 603 820 604 821
rect 605 820 606 821
rect 600 821 606 825
rect 600 825 601 826
rect 602 825 603 826
rect 603 825 604 826
rect 605 825 606 826
rect 480 320 481 321
rect 482 320 483 321
rect 483 320 484 321
rect 485 320 486 321
rect 480 321 486 325
rect 480 325 481 326
rect 482 325 483 326
rect 483 325 484 326
rect 485 325 486 326
rect 740 440 741 441
rect 742 440 743 441
rect 743 440 744 441
rect 745 440 746 441
rect 740 441 746 445
rect 740 445 741 446
rect 742 445 743 446
rect 743 445 744 446
rect 745 445 746 446
rect 480 540 481 541
rect 482 540 483 541
rect 483 540 484 541
rect 485 540 486 541
rect 480 541 486 545
rect 480 545 481 546
rect 482 545 483 546
rect 483 545 484 546
rect 485 545 486 546
rect 540 840 541 841
rect 542 840 543 841
rect 543 840 544 841
rect 545 840 546 841
rect 540 841 546 845
rect 540 845 541 846
rect 542 845 543 846
rect 543 845 544 846
rect 545 845 546 846
rect 440 840 441 841
rect 442 840 443 841
rect 443 840 444 841
rect 445 840 446 841
rect 440 841 446 845
rect 440 845 441 846
rect 442 845 443 846
rect 443 845 444 846
rect 445 845 446 846
rect 460 860 461 861
rect 462 860 463 861
rect 463 860 464 861
rect 465 860 466 861
rect 460 861 466 865
rect 460 865 461 866
rect 462 865 463 866
rect 463 865 464 866
rect 465 865 466 866
rect 300 700 301 701
rect 302 700 303 701
rect 303 700 304 701
rect 305 700 306 701
rect 300 701 306 705
rect 300 705 301 706
rect 302 705 303 706
rect 303 705 304 706
rect 305 705 306 706
rect 460 520 461 521
rect 462 520 463 521
rect 463 520 464 521
rect 465 520 466 521
rect 460 521 466 525
rect 460 525 461 526
rect 462 525 463 526
rect 463 525 464 526
rect 465 525 466 526
rect 420 800 421 801
rect 422 800 423 801
rect 423 800 424 801
rect 425 800 426 801
rect 420 801 426 805
rect 420 805 421 806
rect 422 805 423 806
rect 423 805 424 806
rect 425 805 426 806
rect 520 600 521 601
rect 522 600 523 601
rect 523 600 524 601
rect 525 600 526 601
rect 520 601 526 605
rect 520 605 521 606
rect 522 605 523 606
rect 523 605 524 606
rect 525 605 526 606
rect 760 720 761 721
rect 762 720 763 721
rect 763 720 764 721
rect 765 720 766 721
rect 760 721 766 725
rect 760 725 761 726
rect 762 725 763 726
rect 763 725 764 726
rect 765 725 766 726
rect 340 560 341 561
rect 342 560 343 561
rect 343 560 344 561
rect 345 560 346 561
rect 340 561 346 565
rect 340 565 341 566
rect 342 565 343 566
rect 343 565 344 566
rect 345 565 346 566
rect 500 180 501 181
rect 502 180 503 181
rect 503 180 504 181
rect 505 180 506 181
rect 500 181 506 185
rect 500 185 501 186
rect 502 185 503 186
rect 503 185 504 186
rect 505 185 506 186
rect 440 380 441 381
rect 442 380 443 381
rect 443 380 444 381
rect 445 380 446 381
rect 440 381 446 385
rect 440 385 441 386
rect 442 385 443 386
rect 443 385 444 386
rect 445 385 446 386
rect 280 340 281 341
rect 282 340 283 341
rect 283 340 284 341
rect 285 340 286 341
rect 280 341 286 345
rect 280 345 281 346
rect 282 345 283 346
rect 283 345 284 346
rect 285 345 286 346
rect 220 560 221 561
rect 222 560 223 561
rect 223 560 224 561
rect 225 560 226 561
rect 220 561 226 565
rect 220 565 221 566
rect 222 565 223 566
rect 223 565 224 566
rect 225 565 226 566
rect 840 440 841 441
rect 842 440 843 441
rect 843 440 844 441
rect 845 440 846 441
rect 840 441 846 445
rect 840 445 841 446
rect 842 445 843 446
rect 843 445 844 446
rect 845 445 846 446
rect 240 680 241 681
rect 242 680 243 681
rect 243 680 244 681
rect 245 680 246 681
rect 240 681 246 685
rect 240 685 241 686
rect 242 685 243 686
rect 243 685 244 686
rect 245 685 246 686
rect 500 600 501 601
rect 502 600 503 601
rect 503 600 504 601
rect 505 600 506 601
rect 500 601 506 605
rect 500 605 501 606
rect 502 605 503 606
rect 503 605 504 606
rect 505 605 506 606
rect 740 740 741 741
rect 742 740 743 741
rect 743 740 744 741
rect 745 740 746 741
rect 740 741 746 745
rect 740 745 741 746
rect 742 745 743 746
rect 743 745 744 746
rect 745 745 746 746
rect 200 360 201 361
rect 202 360 203 361
rect 203 360 204 361
rect 205 360 206 361
rect 200 361 206 365
rect 200 365 201 366
rect 202 365 203 366
rect 203 365 204 366
rect 205 365 206 366
rect 160 620 161 621
rect 162 620 163 621
rect 163 620 164 621
rect 165 620 166 621
rect 160 621 166 625
rect 160 625 161 626
rect 162 625 163 626
rect 163 625 164 626
rect 165 625 166 626
rect 280 580 281 581
rect 282 580 283 581
rect 283 580 284 581
rect 285 580 286 581
rect 280 581 286 585
rect 280 585 281 586
rect 282 585 283 586
rect 283 585 284 586
rect 285 585 286 586
rect 740 600 741 601
rect 742 600 743 601
rect 743 600 744 601
rect 745 600 746 601
rect 740 601 746 605
rect 740 605 741 606
rect 742 605 743 606
rect 743 605 744 606
rect 745 605 746 606
rect 460 840 461 841
rect 462 840 463 841
rect 463 840 464 841
rect 465 840 466 841
rect 460 841 466 845
rect 460 845 461 846
rect 462 845 463 846
rect 463 845 464 846
rect 465 845 466 846
rect 680 380 681 381
rect 682 380 683 381
rect 683 380 684 381
rect 685 380 686 381
rect 680 381 686 385
rect 680 385 681 386
rect 682 385 683 386
rect 683 385 684 386
rect 685 385 686 386
rect 240 440 241 441
rect 242 440 243 441
rect 243 440 244 441
rect 245 440 246 441
rect 240 441 246 445
rect 240 445 241 446
rect 242 445 243 446
rect 243 445 244 446
rect 245 445 246 446
rect 640 780 641 781
rect 642 780 643 781
rect 643 780 644 781
rect 645 780 646 781
rect 640 781 646 785
rect 640 785 641 786
rect 642 785 643 786
rect 643 785 644 786
rect 645 785 646 786
rect 460 340 461 341
rect 462 340 463 341
rect 463 340 464 341
rect 465 340 466 341
rect 460 341 466 345
rect 460 345 461 346
rect 462 345 463 346
rect 463 345 464 346
rect 465 345 466 346
rect 740 660 741 661
rect 742 660 743 661
rect 743 660 744 661
rect 745 660 746 661
rect 740 661 746 665
rect 740 665 741 666
rect 742 665 743 666
rect 743 665 744 666
rect 745 665 746 666
rect 360 600 361 601
rect 362 600 363 601
rect 363 600 364 601
rect 365 600 366 601
rect 360 601 366 605
rect 360 605 361 606
rect 362 605 363 606
rect 363 605 364 606
rect 365 605 366 606
rect 420 480 421 481
rect 422 480 423 481
rect 423 480 424 481
rect 425 480 426 481
rect 420 481 426 485
rect 420 485 421 486
rect 422 485 423 486
rect 423 485 424 486
rect 425 485 426 486
rect 700 660 701 661
rect 702 660 703 661
rect 703 660 704 661
rect 705 660 706 661
rect 700 661 706 665
rect 700 665 701 666
rect 702 665 703 666
rect 703 665 704 666
rect 705 665 706 666
rect 340 320 341 321
rect 342 320 343 321
rect 343 320 344 321
rect 345 320 346 321
rect 340 321 346 325
rect 340 325 341 326
rect 342 325 343 326
rect 343 325 344 326
rect 345 325 346 326
rect 540 540 541 541
rect 542 540 543 541
rect 543 540 544 541
rect 545 540 546 541
rect 540 541 546 545
rect 540 545 541 546
rect 542 545 543 546
rect 543 545 544 546
rect 545 545 546 546
rect 220 460 221 461
rect 222 460 223 461
rect 223 460 224 461
rect 225 460 226 461
rect 220 461 226 465
rect 220 465 221 466
rect 222 465 223 466
rect 223 465 224 466
rect 225 465 226 466
rect 860 460 861 461
rect 862 460 863 461
rect 863 460 864 461
rect 865 460 866 461
rect 860 461 866 465
rect 860 465 861 466
rect 862 465 863 466
rect 863 465 864 466
rect 865 465 866 466
rect 560 740 561 741
rect 562 740 563 741
rect 563 740 564 741
rect 565 740 566 741
rect 560 741 566 745
rect 560 745 561 746
rect 562 745 563 746
rect 563 745 564 746
rect 565 745 566 746
rect 160 600 161 601
rect 162 600 163 601
rect 163 600 164 601
rect 165 600 166 601
rect 160 601 166 605
rect 160 605 161 606
rect 162 605 163 606
rect 163 605 164 606
rect 165 605 166 606
rect 640 260 641 261
rect 642 260 643 261
rect 643 260 644 261
rect 645 260 646 261
rect 640 261 646 265
rect 640 265 641 266
rect 642 265 643 266
rect 643 265 644 266
rect 645 265 646 266
rect 720 260 721 261
rect 722 260 723 261
rect 723 260 724 261
rect 725 260 726 261
rect 720 261 726 265
rect 720 265 721 266
rect 722 265 723 266
rect 723 265 724 266
rect 725 265 726 266
rect 780 540 781 541
rect 782 540 783 541
rect 783 540 784 541
rect 785 540 786 541
rect 780 541 786 545
rect 780 545 781 546
rect 782 545 783 546
rect 783 545 784 546
rect 785 545 786 546
rect 560 720 561 721
rect 562 720 563 721
rect 563 720 564 721
rect 565 720 566 721
rect 560 721 566 725
rect 560 725 561 726
rect 562 725 563 726
rect 563 725 564 726
rect 565 725 566 726
rect 500 260 501 261
rect 502 260 503 261
rect 503 260 504 261
rect 505 260 506 261
rect 500 261 506 265
rect 500 265 501 266
rect 502 265 503 266
rect 503 265 504 266
rect 505 265 506 266
rect 240 640 241 641
rect 242 640 243 641
rect 243 640 244 641
rect 245 640 246 641
rect 240 641 246 645
rect 240 645 241 646
rect 242 645 243 646
rect 243 645 244 646
rect 245 645 246 646
rect 460 400 461 401
rect 462 400 463 401
rect 463 400 464 401
rect 465 400 466 401
rect 460 401 466 405
rect 460 405 461 406
rect 462 405 463 406
rect 463 405 464 406
rect 465 405 466 406
rect 740 320 741 321
rect 742 320 743 321
rect 743 320 744 321
rect 745 320 746 321
rect 740 321 746 325
rect 740 325 741 326
rect 742 325 743 326
rect 743 325 744 326
rect 745 325 746 326
rect 360 700 361 701
rect 362 700 363 701
rect 363 700 364 701
rect 365 700 366 701
rect 360 701 366 705
rect 360 705 361 706
rect 362 705 363 706
rect 363 705 364 706
rect 365 705 366 706
rect 440 720 441 721
rect 442 720 443 721
rect 443 720 444 721
rect 445 720 446 721
rect 440 721 446 725
rect 440 725 441 726
rect 442 725 443 726
rect 443 725 444 726
rect 445 725 446 726
rect 400 620 401 621
rect 402 620 403 621
rect 403 620 404 621
rect 405 620 406 621
rect 400 621 406 625
rect 400 625 401 626
rect 402 625 403 626
rect 403 625 404 626
rect 405 625 406 626
rect 420 420 421 421
rect 422 420 423 421
rect 423 420 424 421
rect 425 420 426 421
rect 420 421 426 425
rect 420 425 421 426
rect 422 425 423 426
rect 423 425 424 426
rect 425 425 426 426
rect 220 400 221 401
rect 222 400 223 401
rect 223 400 224 401
rect 225 400 226 401
rect 220 401 226 405
rect 220 405 221 406
rect 222 405 223 406
rect 223 405 224 406
rect 225 405 226 406
rect 740 580 741 581
rect 742 580 743 581
rect 743 580 744 581
rect 745 580 746 581
rect 740 581 746 585
rect 740 585 741 586
rect 742 585 743 586
rect 743 585 744 586
rect 745 585 746 586
rect 460 260 461 261
rect 462 260 463 261
rect 463 260 464 261
rect 465 260 466 261
rect 460 261 466 265
rect 460 265 461 266
rect 462 265 463 266
rect 463 265 464 266
rect 465 265 466 266
rect 740 520 741 521
rect 742 520 743 521
rect 743 520 744 521
rect 745 520 746 521
rect 740 521 746 525
rect 740 525 741 526
rect 742 525 743 526
rect 743 525 744 526
rect 745 525 746 526
rect 460 780 461 781
rect 462 780 463 781
rect 463 780 464 781
rect 465 780 466 781
rect 460 781 466 785
rect 460 785 461 786
rect 462 785 463 786
rect 463 785 464 786
rect 465 785 466 786
rect 100 560 101 561
rect 102 560 103 561
rect 103 560 104 561
rect 105 560 106 561
rect 100 561 106 565
rect 100 565 101 566
rect 102 565 103 566
rect 103 565 104 566
rect 105 565 106 566
rect 480 720 481 721
rect 482 720 483 721
rect 483 720 484 721
rect 485 720 486 721
rect 480 721 486 725
rect 480 725 481 726
rect 482 725 483 726
rect 483 725 484 726
rect 485 725 486 726
rect 580 680 581 681
rect 582 680 583 681
rect 583 680 584 681
rect 585 680 586 681
rect 580 681 586 685
rect 580 685 581 686
rect 582 685 583 686
rect 583 685 584 686
rect 585 685 586 686
rect 540 760 541 761
rect 542 760 543 761
rect 543 760 544 761
rect 545 760 546 761
rect 540 761 546 765
rect 540 765 541 766
rect 542 765 543 766
rect 543 765 544 766
rect 545 765 546 766
rect 420 280 421 281
rect 422 280 423 281
rect 423 280 424 281
rect 425 280 426 281
rect 420 281 426 285
rect 420 285 421 286
rect 422 285 423 286
rect 423 285 424 286
rect 425 285 426 286
rect 680 240 681 241
rect 682 240 683 241
rect 683 240 684 241
rect 685 240 686 241
rect 680 241 686 245
rect 680 245 681 246
rect 682 245 683 246
rect 683 245 684 246
rect 685 245 686 246
rect 160 500 161 501
rect 162 500 163 501
rect 163 500 164 501
rect 165 500 166 501
rect 160 501 166 505
rect 160 505 161 506
rect 162 505 163 506
rect 163 505 164 506
rect 165 505 166 506
rect 640 520 641 521
rect 642 520 643 521
rect 643 520 644 521
rect 645 520 646 521
rect 640 521 646 525
rect 640 525 641 526
rect 642 525 643 526
rect 643 525 644 526
rect 645 525 646 526
rect 860 480 861 481
rect 862 480 863 481
rect 863 480 864 481
rect 865 480 866 481
rect 860 481 866 485
rect 860 485 861 486
rect 862 485 863 486
rect 863 485 864 486
rect 865 485 866 486
rect 680 720 681 721
rect 682 720 683 721
rect 683 720 684 721
rect 685 720 686 721
rect 680 721 686 725
rect 680 725 681 726
rect 682 725 683 726
rect 683 725 684 726
rect 685 725 686 726
rect 460 180 461 181
rect 462 180 463 181
rect 463 180 464 181
rect 465 180 466 181
rect 460 181 466 185
rect 460 185 461 186
rect 462 185 463 186
rect 463 185 464 186
rect 465 185 466 186
rect 560 860 561 861
rect 562 860 563 861
rect 563 860 564 861
rect 565 860 566 861
rect 560 861 566 865
rect 560 865 561 866
rect 562 865 563 866
rect 563 865 564 866
rect 565 865 566 866
rect 240 360 241 361
rect 242 360 243 361
rect 243 360 244 361
rect 245 360 246 361
rect 240 361 246 365
rect 240 365 241 366
rect 242 365 243 366
rect 243 365 244 366
rect 245 365 246 366
rect 700 280 701 281
rect 702 280 703 281
rect 703 280 704 281
rect 705 280 706 281
rect 700 281 706 285
rect 700 285 701 286
rect 702 285 703 286
rect 703 285 704 286
rect 705 285 706 286
rect 260 700 261 701
rect 262 700 263 701
rect 263 700 264 701
rect 265 700 266 701
rect 260 701 266 705
rect 260 705 261 706
rect 262 705 263 706
rect 263 705 264 706
rect 265 705 266 706
rect 140 440 141 441
rect 142 440 143 441
rect 143 440 144 441
rect 145 440 146 441
rect 140 441 146 445
rect 140 445 141 446
rect 142 445 143 446
rect 143 445 144 446
rect 145 445 146 446
rect 240 540 241 541
rect 242 540 243 541
rect 243 540 244 541
rect 245 540 246 541
rect 240 541 246 545
rect 240 545 241 546
rect 242 545 243 546
rect 243 545 244 546
rect 245 545 246 546
rect 840 620 841 621
rect 842 620 843 621
rect 843 620 844 621
rect 845 620 846 621
rect 840 621 846 625
rect 840 625 841 626
rect 842 625 843 626
rect 843 625 844 626
rect 845 625 846 626
rect 780 340 781 341
rect 782 340 783 341
rect 783 340 784 341
rect 785 340 786 341
rect 780 341 786 345
rect 780 345 781 346
rect 782 345 783 346
rect 783 345 784 346
rect 785 345 786 346
rect 220 420 221 421
rect 222 420 223 421
rect 223 420 224 421
rect 225 420 226 421
rect 220 421 226 425
rect 220 425 221 426
rect 222 425 223 426
rect 223 425 224 426
rect 225 425 226 426
rect 560 280 561 281
rect 562 280 563 281
rect 563 280 564 281
rect 565 280 566 281
rect 560 281 566 285
rect 560 285 561 286
rect 562 285 563 286
rect 563 285 564 286
rect 565 285 566 286
rect 460 420 461 421
rect 462 420 463 421
rect 463 420 464 421
rect 465 420 466 421
rect 460 421 466 425
rect 460 425 461 426
rect 462 425 463 426
rect 463 425 464 426
rect 465 425 466 426
rect 420 700 421 701
rect 422 700 423 701
rect 423 700 424 701
rect 425 700 426 701
rect 420 701 426 705
rect 420 705 421 706
rect 422 705 423 706
rect 423 705 424 706
rect 425 705 426 706
rect 140 560 141 561
rect 142 560 143 561
rect 143 560 144 561
rect 145 560 146 561
rect 140 561 146 565
rect 140 565 141 566
rect 142 565 143 566
rect 143 565 144 566
rect 145 565 146 566
rect 680 500 681 501
rect 682 500 683 501
rect 683 500 684 501
rect 685 500 686 501
rect 680 501 686 505
rect 680 505 681 506
rect 682 505 683 506
rect 683 505 684 506
rect 685 505 686 506
rect 820 560 821 561
rect 822 560 823 561
rect 823 560 824 561
rect 825 560 826 561
rect 820 561 826 565
rect 820 565 821 566
rect 822 565 823 566
rect 823 565 824 566
rect 825 565 826 566
rect 560 320 561 321
rect 562 320 563 321
rect 563 320 564 321
rect 565 320 566 321
rect 560 321 566 325
rect 560 325 561 326
rect 562 325 563 326
rect 563 325 564 326
rect 565 325 566 326
rect 840 580 841 581
rect 842 580 843 581
rect 843 580 844 581
rect 845 580 846 581
rect 840 581 846 585
rect 840 585 841 586
rect 842 585 843 586
rect 843 585 844 586
rect 845 585 846 586
rect 560 760 561 761
rect 562 760 563 761
rect 563 760 564 761
rect 565 760 566 761
rect 560 761 566 765
rect 560 765 561 766
rect 562 765 563 766
rect 563 765 564 766
rect 565 765 566 766
rect 700 680 701 681
rect 702 680 703 681
rect 703 680 704 681
rect 705 680 706 681
rect 700 681 706 685
rect 700 685 701 686
rect 702 685 703 686
rect 703 685 704 686
rect 705 685 706 686
rect 440 600 441 601
rect 442 600 443 601
rect 443 600 444 601
rect 445 600 446 601
rect 440 601 446 605
rect 440 605 441 606
rect 442 605 443 606
rect 443 605 444 606
rect 445 605 446 606
rect 500 780 501 781
rect 502 780 503 781
rect 503 780 504 781
rect 505 780 506 781
rect 500 781 506 785
rect 500 785 501 786
rect 502 785 503 786
rect 503 785 504 786
rect 505 785 506 786
rect 500 220 501 221
rect 502 220 503 221
rect 503 220 504 221
rect 505 220 506 221
rect 500 221 506 225
rect 500 225 501 226
rect 502 225 503 226
rect 503 225 504 226
rect 505 225 506 226
rect 260 460 261 461
rect 262 460 263 461
rect 263 460 264 461
rect 265 460 266 461
rect 260 461 266 465
rect 260 465 261 466
rect 262 465 263 466
rect 263 465 264 466
rect 265 465 266 466
rect 540 260 541 261
rect 542 260 543 261
rect 543 260 544 261
rect 545 260 546 261
rect 540 261 546 265
rect 540 265 541 266
rect 542 265 543 266
rect 543 265 544 266
rect 545 265 546 266
rect 660 280 661 281
rect 662 280 663 281
rect 663 280 664 281
rect 665 280 666 281
rect 660 281 666 285
rect 660 285 661 286
rect 662 285 663 286
rect 663 285 664 286
rect 665 285 666 286
rect 620 220 621 221
rect 622 220 623 221
rect 623 220 624 221
rect 625 220 626 221
rect 620 221 626 225
rect 620 225 621 226
rect 622 225 623 226
rect 623 225 624 226
rect 625 225 626 226
rect 720 280 721 281
rect 722 280 723 281
rect 723 280 724 281
rect 725 280 726 281
rect 720 281 726 285
rect 720 285 721 286
rect 722 285 723 286
rect 723 285 724 286
rect 725 285 726 286
rect 680 560 681 561
rect 682 560 683 561
rect 683 560 684 561
rect 685 560 686 561
rect 680 561 686 565
rect 680 565 681 566
rect 682 565 683 566
rect 683 565 684 566
rect 685 565 686 566
rect 700 620 701 621
rect 702 620 703 621
rect 703 620 704 621
rect 705 620 706 621
rect 700 621 706 625
rect 700 625 701 626
rect 702 625 703 626
rect 703 625 704 626
rect 705 625 706 626
rect 820 780 821 781
rect 822 780 823 781
rect 823 780 824 781
rect 825 780 826 781
rect 820 781 826 785
rect 820 785 821 786
rect 822 785 823 786
rect 823 785 824 786
rect 825 785 826 786
rect 240 420 241 421
rect 242 420 243 421
rect 243 420 244 421
rect 245 420 246 421
rect 240 421 246 425
rect 240 425 241 426
rect 242 425 243 426
rect 243 425 244 426
rect 245 425 246 426
rect 340 300 341 301
rect 342 300 343 301
rect 343 300 344 301
rect 345 300 346 301
rect 340 301 346 305
rect 340 305 341 306
rect 342 305 343 306
rect 343 305 344 306
rect 345 305 346 306
rect 580 160 581 161
rect 582 160 583 161
rect 583 160 584 161
rect 585 160 586 161
rect 580 161 586 165
rect 580 165 581 166
rect 582 165 583 166
rect 583 165 584 166
rect 585 165 586 166
rect 500 680 501 681
rect 502 680 503 681
rect 503 680 504 681
rect 505 680 506 681
rect 500 681 506 685
rect 500 685 501 686
rect 502 685 503 686
rect 503 685 504 686
rect 505 685 506 686
rect 820 400 821 401
rect 822 400 823 401
rect 823 400 824 401
rect 825 400 826 401
rect 820 401 826 405
rect 820 405 821 406
rect 822 405 823 406
rect 823 405 824 406
rect 825 405 826 406
rect 420 500 421 501
rect 422 500 423 501
rect 423 500 424 501
rect 425 500 426 501
rect 420 501 426 505
rect 420 505 421 506
rect 422 505 423 506
rect 423 505 424 506
rect 425 505 426 506
rect 700 420 701 421
rect 702 420 703 421
rect 703 420 704 421
rect 705 420 706 421
rect 700 421 706 425
rect 700 425 701 426
rect 702 425 703 426
rect 703 425 704 426
rect 705 425 706 426
rect 620 200 621 201
rect 622 200 623 201
rect 623 200 624 201
rect 625 200 626 201
rect 620 201 626 205
rect 620 205 621 206
rect 622 205 623 206
rect 623 205 624 206
rect 625 205 626 206
rect 480 220 481 221
rect 482 220 483 221
rect 483 220 484 221
rect 485 220 486 221
rect 480 221 486 225
rect 480 225 481 226
rect 482 225 483 226
rect 483 225 484 226
rect 485 225 486 226
rect 140 540 141 541
rect 142 540 143 541
rect 143 540 144 541
rect 145 540 146 541
rect 140 541 146 545
rect 140 545 141 546
rect 142 545 143 546
rect 143 545 144 546
rect 145 545 146 546
rect 240 660 241 661
rect 242 660 243 661
rect 243 660 244 661
rect 245 660 246 661
rect 240 661 246 665
rect 240 665 241 666
rect 242 665 243 666
rect 243 665 244 666
rect 245 665 246 666
rect 540 200 541 201
rect 542 200 543 201
rect 543 200 544 201
rect 545 200 546 201
rect 540 201 546 205
rect 540 205 541 206
rect 542 205 543 206
rect 543 205 544 206
rect 545 205 546 206
rect 380 420 381 421
rect 382 420 383 421
rect 383 420 384 421
rect 385 420 386 421
rect 380 421 386 425
rect 380 425 381 426
rect 382 425 383 426
rect 383 425 384 426
rect 385 425 386 426
rect 440 820 441 821
rect 442 820 443 821
rect 443 820 444 821
rect 445 820 446 821
rect 440 821 446 825
rect 440 825 441 826
rect 442 825 443 826
rect 443 825 444 826
rect 445 825 446 826
rect 280 400 281 401
rect 282 400 283 401
rect 283 400 284 401
rect 285 400 286 401
rect 280 401 286 405
rect 280 405 281 406
rect 282 405 283 406
rect 283 405 284 406
rect 285 405 286 406
rect 660 240 661 241
rect 662 240 663 241
rect 663 240 664 241
rect 665 240 666 241
rect 660 241 666 245
rect 660 245 661 246
rect 662 245 663 246
rect 663 245 664 246
rect 665 245 666 246
rect 220 600 221 601
rect 222 600 223 601
rect 223 600 224 601
rect 225 600 226 601
rect 220 601 226 605
rect 220 605 221 606
rect 222 605 223 606
rect 223 605 224 606
rect 225 605 226 606
rect 460 300 461 301
rect 462 300 463 301
rect 463 300 464 301
rect 465 300 466 301
rect 460 301 466 305
rect 460 305 461 306
rect 462 305 463 306
rect 463 305 464 306
rect 465 305 466 306
rect 180 420 181 421
rect 182 420 183 421
rect 183 420 184 421
rect 185 420 186 421
rect 180 421 186 425
rect 180 425 181 426
rect 182 425 183 426
rect 183 425 184 426
rect 185 425 186 426
rect 380 260 381 261
rect 382 260 383 261
rect 383 260 384 261
rect 385 260 386 261
rect 380 261 386 265
rect 380 265 381 266
rect 382 265 383 266
rect 383 265 384 266
rect 385 265 386 266
rect 300 320 301 321
rect 302 320 303 321
rect 303 320 304 321
rect 305 320 306 321
rect 300 321 306 325
rect 300 325 301 326
rect 302 325 303 326
rect 303 325 304 326
rect 305 325 306 326
rect 180 560 181 561
rect 182 560 183 561
rect 183 560 184 561
rect 185 560 186 561
rect 180 561 186 565
rect 180 565 181 566
rect 182 565 183 566
rect 183 565 184 566
rect 185 565 186 566
rect 380 680 381 681
rect 382 680 383 681
rect 383 680 384 681
rect 385 680 386 681
rect 380 681 386 685
rect 380 685 381 686
rect 382 685 383 686
rect 383 685 384 686
rect 385 685 386 686
rect 840 500 841 501
rect 842 500 843 501
rect 843 500 844 501
rect 845 500 846 501
rect 840 501 846 505
rect 840 505 841 506
rect 842 505 843 506
rect 843 505 844 506
rect 845 505 846 506
rect 460 640 461 641
rect 462 640 463 641
rect 463 640 464 641
rect 465 640 466 641
rect 460 641 466 645
rect 460 645 461 646
rect 462 645 463 646
rect 463 645 464 646
rect 465 645 466 646
rect 520 640 521 641
rect 522 640 523 641
rect 523 640 524 641
rect 525 640 526 641
rect 520 641 526 645
rect 520 645 521 646
rect 522 645 523 646
rect 523 645 524 646
rect 525 645 526 646
rect 760 360 761 361
rect 762 360 763 361
rect 763 360 764 361
rect 765 360 766 361
rect 760 361 766 365
rect 760 365 761 366
rect 762 365 763 366
rect 763 365 764 366
rect 765 365 766 366
rect 340 780 341 781
rect 342 780 343 781
rect 343 780 344 781
rect 345 780 346 781
rect 340 781 346 785
rect 340 785 341 786
rect 342 785 343 786
rect 343 785 344 786
rect 345 785 346 786
rect 620 440 621 441
rect 622 440 623 441
rect 623 440 624 441
rect 625 440 626 441
rect 620 441 626 445
rect 620 445 621 446
rect 622 445 623 446
rect 623 445 624 446
rect 625 445 626 446
rect 520 280 521 281
rect 522 280 523 281
rect 523 280 524 281
rect 525 280 526 281
rect 520 281 526 285
rect 520 285 521 286
rect 522 285 523 286
rect 523 285 524 286
rect 525 285 526 286
rect 500 400 501 401
rect 502 400 503 401
rect 503 400 504 401
rect 505 400 506 401
rect 500 401 506 405
rect 500 405 501 406
rect 502 405 503 406
rect 503 405 504 406
rect 505 405 506 406
rect 340 580 341 581
rect 342 580 343 581
rect 343 580 344 581
rect 345 580 346 581
rect 340 581 346 585
rect 340 585 341 586
rect 342 585 343 586
rect 343 585 344 586
rect 345 585 346 586
rect 820 480 821 481
rect 822 480 823 481
rect 823 480 824 481
rect 825 480 826 481
rect 820 481 826 485
rect 820 485 821 486
rect 822 485 823 486
rect 823 485 824 486
rect 825 485 826 486
rect 540 480 541 481
rect 542 480 543 481
rect 543 480 544 481
rect 545 480 546 481
rect 540 481 546 485
rect 540 485 541 486
rect 542 485 543 486
rect 543 485 544 486
rect 545 485 546 486
rect 340 380 341 381
rect 342 380 343 381
rect 343 380 344 381
rect 345 380 346 381
rect 340 381 346 385
rect 340 385 341 386
rect 342 385 343 386
rect 343 385 344 386
rect 345 385 346 386
rect 460 460 461 461
rect 462 460 463 461
rect 463 460 464 461
rect 465 460 466 461
rect 460 461 466 465
rect 460 465 461 466
rect 462 465 463 466
rect 463 465 464 466
rect 465 465 466 466
rect 560 240 561 241
rect 562 240 563 241
rect 563 240 564 241
rect 565 240 566 241
rect 560 241 566 245
rect 560 245 561 246
rect 562 245 563 246
rect 563 245 564 246
rect 565 245 566 246
rect 600 780 601 781
rect 602 780 603 781
rect 603 780 604 781
rect 605 780 606 781
rect 600 781 606 785
rect 600 785 601 786
rect 602 785 603 786
rect 603 785 604 786
rect 605 785 606 786
rect 500 660 501 661
rect 502 660 503 661
rect 503 660 504 661
rect 505 660 506 661
rect 500 661 506 665
rect 500 665 501 666
rect 502 665 503 666
rect 503 665 504 666
rect 505 665 506 666
rect 280 480 281 481
rect 282 480 283 481
rect 283 480 284 481
rect 285 480 286 481
rect 280 481 286 485
rect 280 485 281 486
rect 282 485 283 486
rect 283 485 284 486
rect 285 485 286 486
rect 780 440 781 441
rect 782 440 783 441
rect 783 440 784 441
rect 785 440 786 441
rect 780 441 786 445
rect 780 445 781 446
rect 782 445 783 446
rect 783 445 784 446
rect 785 445 786 446
rect 480 240 481 241
rect 482 240 483 241
rect 483 240 484 241
rect 485 240 486 241
rect 480 241 486 245
rect 480 245 481 246
rect 482 245 483 246
rect 483 245 484 246
rect 485 245 486 246
rect 700 740 701 741
rect 702 740 703 741
rect 703 740 704 741
rect 705 740 706 741
rect 700 741 706 745
rect 700 745 701 746
rect 702 745 703 746
rect 703 745 704 746
rect 705 745 706 746
rect 540 400 541 401
rect 542 400 543 401
rect 543 400 544 401
rect 545 400 546 401
rect 540 401 546 405
rect 540 405 541 406
rect 542 405 543 406
rect 543 405 544 406
rect 545 405 546 406
rect 440 160 441 161
rect 442 160 443 161
rect 443 160 444 161
rect 445 160 446 161
rect 440 161 446 165
rect 440 165 441 166
rect 442 165 443 166
rect 443 165 444 166
rect 445 165 446 166
rect 120 600 121 601
rect 122 600 123 601
rect 123 600 124 601
rect 125 600 126 601
rect 120 601 126 605
rect 120 605 121 606
rect 122 605 123 606
rect 123 605 124 606
rect 125 605 126 606
rect 700 580 701 581
rect 702 580 703 581
rect 703 580 704 581
rect 705 580 706 581
rect 700 581 706 585
rect 700 585 701 586
rect 702 585 703 586
rect 703 585 704 586
rect 705 585 706 586
rect 460 540 461 541
rect 462 540 463 541
rect 463 540 464 541
rect 465 540 466 541
rect 460 541 466 545
rect 460 545 461 546
rect 462 545 463 546
rect 463 545 464 546
rect 465 545 466 546
rect 400 300 401 301
rect 402 300 403 301
rect 403 300 404 301
rect 405 300 406 301
rect 400 301 406 305
rect 400 305 401 306
rect 402 305 403 306
rect 403 305 404 306
rect 405 305 406 306
rect 320 320 321 321
rect 322 320 323 321
rect 323 320 324 321
rect 325 320 326 321
rect 320 321 326 325
rect 320 325 321 326
rect 322 325 323 326
rect 323 325 324 326
rect 325 325 326 326
rect 260 580 261 581
rect 262 580 263 581
rect 263 580 264 581
rect 265 580 266 581
rect 260 581 266 585
rect 260 585 261 586
rect 262 585 263 586
rect 263 585 264 586
rect 265 585 266 586
rect 560 600 561 601
rect 562 600 563 601
rect 563 600 564 601
rect 565 600 566 601
rect 560 601 566 605
rect 560 605 561 606
rect 562 605 563 606
rect 563 605 564 606
rect 565 605 566 606
rect 640 180 641 181
rect 642 180 643 181
rect 643 180 644 181
rect 645 180 646 181
rect 640 181 646 185
rect 640 185 641 186
rect 642 185 643 186
rect 643 185 644 186
rect 645 185 646 186
rect 720 760 721 761
rect 722 760 723 761
rect 723 760 724 761
rect 725 760 726 761
rect 720 761 726 765
rect 720 765 721 766
rect 722 765 723 766
rect 723 765 724 766
rect 725 765 726 766
rect 120 460 121 461
rect 122 460 123 461
rect 123 460 124 461
rect 125 460 126 461
rect 120 461 126 465
rect 120 465 121 466
rect 122 465 123 466
rect 123 465 124 466
rect 125 465 126 466
rect 400 600 401 601
rect 402 600 403 601
rect 403 600 404 601
rect 405 600 406 601
rect 400 601 406 605
rect 400 605 401 606
rect 402 605 403 606
rect 403 605 404 606
rect 405 605 406 606
rect 520 400 521 401
rect 522 400 523 401
rect 523 400 524 401
rect 525 400 526 401
rect 520 401 526 405
rect 520 405 521 406
rect 522 405 523 406
rect 523 405 524 406
rect 525 405 526 406
rect 680 200 681 201
rect 682 200 683 201
rect 683 200 684 201
rect 685 200 686 201
rect 680 201 686 205
rect 680 205 681 206
rect 682 205 683 206
rect 683 205 684 206
rect 685 205 686 206
rect 620 520 621 521
rect 622 520 623 521
rect 623 520 624 521
rect 625 520 626 521
rect 620 521 626 525
rect 620 525 621 526
rect 622 525 623 526
rect 623 525 624 526
rect 625 525 626 526
rect 260 600 261 601
rect 262 600 263 601
rect 263 600 264 601
rect 265 600 266 601
rect 260 601 266 605
rect 260 605 261 606
rect 262 605 263 606
rect 263 605 264 606
rect 265 605 266 606
rect 520 740 521 741
rect 522 740 523 741
rect 523 740 524 741
rect 525 740 526 741
rect 520 741 526 745
rect 520 745 521 746
rect 522 745 523 746
rect 523 745 524 746
rect 525 745 526 746
rect 620 420 621 421
rect 622 420 623 421
rect 623 420 624 421
rect 625 420 626 421
rect 620 421 626 425
rect 620 425 621 426
rect 622 425 623 426
rect 623 425 624 426
rect 625 425 626 426
rect 280 680 281 681
rect 282 680 283 681
rect 283 680 284 681
rect 285 680 286 681
rect 280 681 286 685
rect 280 685 281 686
rect 282 685 283 686
rect 283 685 284 686
rect 285 685 286 686
rect 420 640 421 641
rect 422 640 423 641
rect 423 640 424 641
rect 425 640 426 641
rect 420 641 426 645
rect 420 645 421 646
rect 422 645 423 646
rect 423 645 424 646
rect 425 645 426 646
rect 560 300 561 301
rect 562 300 563 301
rect 563 300 564 301
rect 565 300 566 301
rect 560 301 566 305
rect 560 305 561 306
rect 562 305 563 306
rect 563 305 564 306
rect 565 305 566 306
rect 320 680 321 681
rect 322 680 323 681
rect 323 680 324 681
rect 325 680 326 681
rect 320 681 326 685
rect 320 685 321 686
rect 322 685 323 686
rect 323 685 324 686
rect 325 685 326 686
rect 560 500 561 501
rect 562 500 563 501
rect 563 500 564 501
rect 565 500 566 501
rect 560 501 566 505
rect 560 505 561 506
rect 562 505 563 506
rect 563 505 564 506
rect 565 505 566 506
rect 240 480 241 481
rect 242 480 243 481
rect 243 480 244 481
rect 245 480 246 481
rect 240 481 246 485
rect 240 485 241 486
rect 242 485 243 486
rect 243 485 244 486
rect 245 485 246 486
rect 700 600 701 601
rect 702 600 703 601
rect 703 600 704 601
rect 705 600 706 601
rect 700 601 706 605
rect 700 605 701 606
rect 702 605 703 606
rect 703 605 704 606
rect 705 605 706 606
rect 280 640 281 641
rect 282 640 283 641
rect 283 640 284 641
rect 285 640 286 641
rect 280 641 286 645
rect 280 645 281 646
rect 282 645 283 646
rect 283 645 284 646
rect 285 645 286 646
rect 300 560 301 561
rect 302 560 303 561
rect 303 560 304 561
rect 305 560 306 561
rect 300 561 306 565
rect 300 565 301 566
rect 302 565 303 566
rect 303 565 304 566
rect 305 565 306 566
rect 440 440 441 441
rect 442 440 443 441
rect 443 440 444 441
rect 445 440 446 441
rect 440 441 446 445
rect 440 445 441 446
rect 442 445 443 446
rect 443 445 444 446
rect 445 445 446 446
rect 600 440 601 441
rect 602 440 603 441
rect 603 440 604 441
rect 605 440 606 441
rect 600 441 606 445
rect 600 445 601 446
rect 602 445 603 446
rect 603 445 604 446
rect 605 445 606 446
rect 620 460 621 461
rect 622 460 623 461
rect 623 460 624 461
rect 625 460 626 461
rect 620 461 626 465
rect 620 465 621 466
rect 622 465 623 466
rect 623 465 624 466
rect 625 465 626 466
rect 660 580 661 581
rect 662 580 663 581
rect 663 580 664 581
rect 665 580 666 581
rect 660 581 666 585
rect 660 585 661 586
rect 662 585 663 586
rect 663 585 664 586
rect 665 585 666 586
rect 400 640 401 641
rect 402 640 403 641
rect 403 640 404 641
rect 405 640 406 641
rect 400 641 406 645
rect 400 645 401 646
rect 402 645 403 646
rect 403 645 404 646
rect 405 645 406 646
rect 260 440 261 441
rect 262 440 263 441
rect 263 440 264 441
rect 265 440 266 441
rect 260 441 266 445
rect 260 445 261 446
rect 262 445 263 446
rect 263 445 264 446
rect 265 445 266 446
rect 860 580 861 581
rect 862 580 863 581
rect 863 580 864 581
rect 865 580 866 581
rect 860 581 866 585
rect 860 585 861 586
rect 862 585 863 586
rect 863 585 864 586
rect 865 585 866 586
rect 720 640 721 641
rect 722 640 723 641
rect 723 640 724 641
rect 725 640 726 641
rect 720 641 726 645
rect 720 645 721 646
rect 722 645 723 646
rect 723 645 724 646
rect 725 645 726 646
rect 380 300 381 301
rect 382 300 383 301
rect 383 300 384 301
rect 385 300 386 301
rect 380 301 386 305
rect 380 305 381 306
rect 382 305 383 306
rect 383 305 384 306
rect 385 305 386 306
rect 420 720 421 721
rect 422 720 423 721
rect 423 720 424 721
rect 425 720 426 721
rect 420 721 426 725
rect 420 725 421 726
rect 422 725 423 726
rect 423 725 424 726
rect 425 725 426 726
rect 300 680 301 681
rect 302 680 303 681
rect 303 680 304 681
rect 305 680 306 681
rect 300 681 306 685
rect 300 685 301 686
rect 302 685 303 686
rect 303 685 304 686
rect 305 685 306 686
rect 620 660 621 661
rect 622 660 623 661
rect 623 660 624 661
rect 625 660 626 661
rect 620 661 626 665
rect 620 665 621 666
rect 622 665 623 666
rect 623 665 624 666
rect 625 665 626 666
rect 700 520 701 521
rect 702 520 703 521
rect 703 520 704 521
rect 705 520 706 521
rect 700 521 706 525
rect 700 525 701 526
rect 702 525 703 526
rect 703 525 704 526
rect 705 525 706 526
rect 320 760 321 761
rect 322 760 323 761
rect 323 760 324 761
rect 325 760 326 761
rect 320 761 326 765
rect 320 765 321 766
rect 322 765 323 766
rect 323 765 324 766
rect 325 765 326 766
rect 480 780 481 781
rect 482 780 483 781
rect 483 780 484 781
rect 485 780 486 781
rect 480 781 486 785
rect 480 785 481 786
rect 482 785 483 786
rect 483 785 484 786
rect 485 785 486 786
rect 700 640 701 641
rect 702 640 703 641
rect 703 640 704 641
rect 705 640 706 641
rect 700 641 706 645
rect 700 645 701 646
rect 702 645 703 646
rect 703 645 704 646
rect 705 645 706 646
rect 580 520 581 521
rect 582 520 583 521
rect 583 520 584 521
rect 585 520 586 521
rect 580 521 586 525
rect 580 525 581 526
rect 582 525 583 526
rect 583 525 584 526
rect 585 525 586 526
rect 600 520 601 521
rect 602 520 603 521
rect 603 520 604 521
rect 605 520 606 521
rect 600 521 606 525
rect 600 525 601 526
rect 602 525 603 526
rect 603 525 604 526
rect 605 525 606 526
rect 460 480 461 481
rect 462 480 463 481
rect 463 480 464 481
rect 465 480 466 481
rect 460 481 466 485
rect 460 485 461 486
rect 462 485 463 486
rect 463 485 464 486
rect 465 485 466 486
rect 600 680 601 681
rect 602 680 603 681
rect 603 680 604 681
rect 605 680 606 681
rect 600 681 606 685
rect 600 685 601 686
rect 602 685 603 686
rect 603 685 604 686
rect 605 685 606 686
rect 480 700 481 701
rect 482 700 483 701
rect 483 700 484 701
rect 485 700 486 701
rect 480 701 486 705
rect 480 705 481 706
rect 482 705 483 706
rect 483 705 484 706
rect 485 705 486 706
rect 760 640 761 641
rect 762 640 763 641
rect 763 640 764 641
rect 765 640 766 641
rect 760 641 766 645
rect 760 645 761 646
rect 762 645 763 646
rect 763 645 764 646
rect 765 645 766 646
rect 420 740 421 741
rect 422 740 423 741
rect 423 740 424 741
rect 425 740 426 741
rect 420 741 426 745
rect 420 745 421 746
rect 422 745 423 746
rect 423 745 424 746
rect 425 745 426 746
rect 700 260 701 261
rect 702 260 703 261
rect 703 260 704 261
rect 705 260 706 261
rect 700 261 706 265
rect 700 265 701 266
rect 702 265 703 266
rect 703 265 704 266
rect 705 265 706 266
rect 440 740 441 741
rect 442 740 443 741
rect 443 740 444 741
rect 445 740 446 741
rect 440 741 446 745
rect 440 745 441 746
rect 442 745 443 746
rect 443 745 444 746
rect 445 745 446 746
rect 380 360 381 361
rect 382 360 383 361
rect 383 360 384 361
rect 385 360 386 361
rect 380 361 386 365
rect 380 365 381 366
rect 382 365 383 366
rect 383 365 384 366
rect 385 365 386 366
rect 340 600 341 601
rect 342 600 343 601
rect 343 600 344 601
rect 345 600 346 601
rect 340 601 346 605
rect 340 605 341 606
rect 342 605 343 606
rect 343 605 344 606
rect 345 605 346 606
rect 560 620 561 621
rect 562 620 563 621
rect 563 620 564 621
rect 565 620 566 621
rect 560 621 566 625
rect 560 625 561 626
rect 562 625 563 626
rect 563 625 564 626
rect 565 625 566 626
rect 640 440 641 441
rect 642 440 643 441
rect 643 440 644 441
rect 645 440 646 441
rect 640 441 646 445
rect 640 445 641 446
rect 642 445 643 446
rect 643 445 644 446
rect 645 445 646 446
rect 320 280 321 281
rect 322 280 323 281
rect 323 280 324 281
rect 325 280 326 281
rect 320 281 326 285
rect 320 285 321 286
rect 322 285 323 286
rect 323 285 324 286
rect 325 285 326 286
rect 660 360 661 361
rect 662 360 663 361
rect 663 360 664 361
rect 665 360 666 361
rect 660 361 666 365
rect 660 365 661 366
rect 662 365 663 366
rect 663 365 664 366
rect 665 365 666 366
rect 300 540 301 541
rect 302 540 303 541
rect 303 540 304 541
rect 305 540 306 541
rect 300 541 306 545
rect 300 545 301 546
rect 302 545 303 546
rect 303 545 304 546
rect 305 545 306 546
rect 400 700 401 701
rect 402 700 403 701
rect 403 700 404 701
rect 405 700 406 701
rect 400 701 406 705
rect 400 705 401 706
rect 402 705 403 706
rect 403 705 404 706
rect 405 705 406 706
rect 620 480 621 481
rect 622 480 623 481
rect 623 480 624 481
rect 625 480 626 481
rect 620 481 626 485
rect 620 485 621 486
rect 622 485 623 486
rect 623 485 624 486
rect 625 485 626 486
rect 540 220 541 221
rect 542 220 543 221
rect 543 220 544 221
rect 545 220 546 221
rect 540 221 546 225
rect 540 225 541 226
rect 542 225 543 226
rect 543 225 544 226
rect 545 225 546 226
rect 580 340 581 341
rect 582 340 583 341
rect 583 340 584 341
rect 585 340 586 341
rect 580 341 586 345
rect 580 345 581 346
rect 582 345 583 346
rect 583 345 584 346
rect 585 345 586 346
rect 500 700 501 701
rect 502 700 503 701
rect 503 700 504 701
rect 505 700 506 701
rect 500 701 506 705
rect 500 705 501 706
rect 502 705 503 706
rect 503 705 504 706
rect 505 705 506 706
rect 480 440 481 441
rect 482 440 483 441
rect 483 440 484 441
rect 485 440 486 441
rect 480 441 486 445
rect 480 445 481 446
rect 482 445 483 446
rect 483 445 484 446
rect 485 445 486 446
rect 720 540 721 541
rect 722 540 723 541
rect 723 540 724 541
rect 725 540 726 541
rect 720 541 726 545
rect 720 545 721 546
rect 722 545 723 546
rect 723 545 724 546
rect 725 545 726 546
rect 300 620 301 621
rect 302 620 303 621
rect 303 620 304 621
rect 305 620 306 621
rect 300 621 306 625
rect 300 625 301 626
rect 302 625 303 626
rect 303 625 304 626
rect 305 625 306 626
rect 860 600 861 601
rect 862 600 863 601
rect 863 600 864 601
rect 865 600 866 601
rect 860 601 866 605
rect 860 605 861 606
rect 862 605 863 606
rect 863 605 864 606
rect 865 605 866 606
rect 520 680 521 681
rect 522 680 523 681
rect 523 680 524 681
rect 525 680 526 681
rect 520 681 526 685
rect 520 685 521 686
rect 522 685 523 686
rect 523 685 524 686
rect 525 685 526 686
rect 760 540 761 541
rect 762 540 763 541
rect 763 540 764 541
rect 765 540 766 541
rect 760 541 766 545
rect 760 545 761 546
rect 762 545 763 546
rect 763 545 764 546
rect 765 545 766 546
rect 220 640 221 641
rect 222 640 223 641
rect 223 640 224 641
rect 225 640 226 641
rect 220 641 226 645
rect 220 645 221 646
rect 222 645 223 646
rect 223 645 224 646
rect 225 645 226 646
rect 300 500 301 501
rect 302 500 303 501
rect 303 500 304 501
rect 305 500 306 501
rect 300 501 306 505
rect 300 505 301 506
rect 302 505 303 506
rect 303 505 304 506
rect 305 505 306 506
rect 400 280 401 281
rect 402 280 403 281
rect 403 280 404 281
rect 405 280 406 281
rect 400 281 406 285
rect 400 285 401 286
rect 402 285 403 286
rect 403 285 404 286
rect 405 285 406 286
rect 440 660 441 661
rect 442 660 443 661
rect 443 660 444 661
rect 445 660 446 661
rect 440 661 446 665
rect 440 665 441 666
rect 442 665 443 666
rect 443 665 444 666
rect 445 665 446 666
rect 540 600 541 601
rect 542 600 543 601
rect 543 600 544 601
rect 545 600 546 601
rect 540 601 546 605
rect 540 605 541 606
rect 542 605 543 606
rect 543 605 544 606
rect 545 605 546 606
rect 360 540 361 541
rect 362 540 363 541
rect 363 540 364 541
rect 365 540 366 541
rect 360 541 366 545
rect 360 545 361 546
rect 362 545 363 546
rect 363 545 364 546
rect 365 545 366 546
rect 340 800 341 801
rect 342 800 343 801
rect 343 800 344 801
rect 345 800 346 801
rect 340 801 346 805
rect 340 805 341 806
rect 342 805 343 806
rect 343 805 344 806
rect 345 805 346 806
rect 580 640 581 641
rect 582 640 583 641
rect 583 640 584 641
rect 585 640 586 641
rect 580 641 586 645
rect 580 645 581 646
rect 582 645 583 646
rect 583 645 584 646
rect 585 645 586 646
rect 500 340 501 341
rect 502 340 503 341
rect 503 340 504 341
rect 505 340 506 341
rect 500 341 506 345
rect 500 345 501 346
rect 502 345 503 346
rect 503 345 504 346
rect 505 345 506 346
rect 200 640 201 641
rect 202 640 203 641
rect 203 640 204 641
rect 205 640 206 641
rect 200 641 206 645
rect 200 645 201 646
rect 202 645 203 646
rect 203 645 204 646
rect 205 645 206 646
rect 660 800 661 801
rect 662 800 663 801
rect 663 800 664 801
rect 665 800 666 801
rect 660 801 666 805
rect 660 805 661 806
rect 662 805 663 806
rect 663 805 664 806
rect 665 805 666 806
rect 160 480 161 481
rect 162 480 163 481
rect 163 480 164 481
rect 165 480 166 481
rect 160 481 166 485
rect 160 485 161 486
rect 162 485 163 486
rect 163 485 164 486
rect 165 485 166 486
rect 300 360 301 361
rect 302 360 303 361
rect 303 360 304 361
rect 305 360 306 361
rect 300 361 306 365
rect 300 365 301 366
rect 302 365 303 366
rect 303 365 304 366
rect 305 365 306 366
rect 420 540 421 541
rect 422 540 423 541
rect 423 540 424 541
rect 425 540 426 541
rect 420 541 426 545
rect 420 545 421 546
rect 422 545 423 546
rect 423 545 424 546
rect 425 545 426 546
rect 620 540 621 541
rect 622 540 623 541
rect 623 540 624 541
rect 625 540 626 541
rect 620 541 626 545
rect 620 545 621 546
rect 622 545 623 546
rect 623 545 624 546
rect 625 545 626 546
rect 460 320 461 321
rect 462 320 463 321
rect 463 320 464 321
rect 465 320 466 321
rect 460 321 466 325
rect 460 325 461 326
rect 462 325 463 326
rect 463 325 464 326
rect 465 325 466 326
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect 520 300 521 301
rect 522 300 523 301
rect 523 300 524 301
rect 525 300 526 301
rect 520 301 526 305
rect 520 305 521 306
rect 522 305 523 306
rect 523 305 524 306
rect 525 305 526 306
rect 640 360 641 361
rect 642 360 643 361
rect 643 360 644 361
rect 645 360 646 361
rect 640 361 646 365
rect 640 365 641 366
rect 642 365 643 366
rect 643 365 644 366
rect 645 365 646 366
rect 220 540 221 541
rect 222 540 223 541
rect 223 540 224 541
rect 225 540 226 541
rect 220 541 226 545
rect 220 545 221 546
rect 222 545 223 546
rect 223 545 224 546
rect 225 545 226 546
rect 400 460 401 461
rect 402 460 403 461
rect 403 460 404 461
rect 405 460 406 461
rect 400 461 406 465
rect 400 465 401 466
rect 402 465 403 466
rect 403 465 404 466
rect 405 465 406 466
rect 640 600 641 601
rect 642 600 643 601
rect 643 600 644 601
rect 645 600 646 601
rect 640 601 646 605
rect 640 605 641 606
rect 642 605 643 606
rect 643 605 644 606
rect 645 605 646 606
rect 880 560 881 561
rect 882 560 883 561
rect 883 560 884 561
rect 885 560 886 561
rect 880 561 886 565
rect 880 565 881 566
rect 882 565 883 566
rect 883 565 884 566
rect 885 565 886 566
rect 340 340 341 341
rect 342 340 343 341
rect 343 340 344 341
rect 345 340 346 341
rect 340 341 346 345
rect 340 345 341 346
rect 342 345 343 346
rect 343 345 344 346
rect 345 345 346 346
rect 700 440 701 441
rect 702 440 703 441
rect 703 440 704 441
rect 705 440 706 441
rect 700 441 706 445
rect 700 445 701 446
rect 702 445 703 446
rect 703 445 704 446
rect 705 445 706 446
rect 420 780 421 781
rect 422 780 423 781
rect 423 780 424 781
rect 425 780 426 781
rect 420 781 426 785
rect 420 785 421 786
rect 422 785 423 786
rect 423 785 424 786
rect 425 785 426 786
rect 360 300 361 301
rect 362 300 363 301
rect 363 300 364 301
rect 365 300 366 301
rect 360 301 366 305
rect 360 305 361 306
rect 362 305 363 306
rect 363 305 364 306
rect 365 305 366 306
rect 540 620 541 621
rect 542 620 543 621
rect 543 620 544 621
rect 545 620 546 621
rect 540 621 546 625
rect 540 625 541 626
rect 542 625 543 626
rect 543 625 544 626
rect 545 625 546 626
rect 360 400 361 401
rect 362 400 363 401
rect 363 400 364 401
rect 365 400 366 401
rect 360 401 366 405
rect 360 405 361 406
rect 362 405 363 406
rect 363 405 364 406
rect 365 405 366 406
rect 260 620 261 621
rect 262 620 263 621
rect 263 620 264 621
rect 265 620 266 621
rect 260 621 266 625
rect 260 625 261 626
rect 262 625 263 626
rect 263 625 264 626
rect 265 625 266 626
rect 640 480 641 481
rect 642 480 643 481
rect 643 480 644 481
rect 645 480 646 481
rect 640 481 646 485
rect 640 485 641 486
rect 642 485 643 486
rect 643 485 644 486
rect 645 485 646 486
rect 640 640 641 641
rect 642 640 643 641
rect 643 640 644 641
rect 645 640 646 641
rect 640 641 646 645
rect 640 645 641 646
rect 642 645 643 646
rect 643 645 644 646
rect 645 645 646 646
rect 400 500 401 501
rect 402 500 403 501
rect 403 500 404 501
rect 405 500 406 501
rect 400 501 406 505
rect 400 505 401 506
rect 402 505 403 506
rect 403 505 404 506
rect 405 505 406 506
rect 580 740 581 741
rect 582 740 583 741
rect 583 740 584 741
rect 585 740 586 741
rect 580 741 586 745
rect 580 745 581 746
rect 582 745 583 746
rect 583 745 584 746
rect 585 745 586 746
rect 140 480 141 481
rect 142 480 143 481
rect 143 480 144 481
rect 145 480 146 481
rect 140 481 146 485
rect 140 485 141 486
rect 142 485 143 486
rect 143 485 144 486
rect 145 485 146 486
rect 660 740 661 741
rect 662 740 663 741
rect 663 740 664 741
rect 665 740 666 741
rect 660 741 666 745
rect 660 745 661 746
rect 662 745 663 746
rect 663 745 664 746
rect 665 745 666 746
rect 400 840 401 841
rect 402 840 403 841
rect 403 840 404 841
rect 405 840 406 841
rect 400 841 406 845
rect 400 845 401 846
rect 402 845 403 846
rect 403 845 404 846
rect 405 845 406 846
rect 380 220 381 221
rect 382 220 383 221
rect 383 220 384 221
rect 385 220 386 221
rect 380 221 386 225
rect 380 225 381 226
rect 382 225 383 226
rect 383 225 384 226
rect 385 225 386 226
rect 340 640 341 641
rect 342 640 343 641
rect 343 640 344 641
rect 345 640 346 641
rect 340 641 346 645
rect 340 645 341 646
rect 342 645 343 646
rect 343 645 344 646
rect 345 645 346 646
rect 200 420 201 421
rect 202 420 203 421
rect 203 420 204 421
rect 205 420 206 421
rect 200 421 206 425
rect 200 425 201 426
rect 202 425 203 426
rect 203 425 204 426
rect 205 425 206 426
rect 760 560 761 561
rect 762 560 763 561
rect 763 560 764 561
rect 765 560 766 561
rect 760 561 766 565
rect 760 565 761 566
rect 762 565 763 566
rect 763 565 764 566
rect 765 565 766 566
rect 300 280 301 281
rect 302 280 303 281
rect 303 280 304 281
rect 305 280 306 281
rect 300 281 306 285
rect 300 285 301 286
rect 302 285 303 286
rect 303 285 304 286
rect 305 285 306 286
rect 180 620 181 621
rect 182 620 183 621
rect 183 620 184 621
rect 185 620 186 621
rect 180 621 186 625
rect 180 625 181 626
rect 182 625 183 626
rect 183 625 184 626
rect 185 625 186 626
rect 420 520 421 521
rect 422 520 423 521
rect 423 520 424 521
rect 425 520 426 521
rect 420 521 426 525
rect 420 525 421 526
rect 422 525 423 526
rect 423 525 424 526
rect 425 525 426 526
rect 540 340 541 341
rect 542 340 543 341
rect 543 340 544 341
rect 545 340 546 341
rect 540 341 546 345
rect 540 345 541 346
rect 542 345 543 346
rect 543 345 544 346
rect 545 345 546 346
rect 640 380 641 381
rect 642 380 643 381
rect 643 380 644 381
rect 645 380 646 381
rect 640 381 646 385
rect 640 385 641 386
rect 642 385 643 386
rect 643 385 644 386
rect 645 385 646 386
rect 800 580 801 581
rect 802 580 803 581
rect 803 580 804 581
rect 805 580 806 581
rect 800 581 806 585
rect 800 585 801 586
rect 802 585 803 586
rect 803 585 804 586
rect 805 585 806 586
rect 240 600 241 601
rect 242 600 243 601
rect 243 600 244 601
rect 245 600 246 601
rect 240 601 246 605
rect 240 605 241 606
rect 242 605 243 606
rect 243 605 244 606
rect 245 605 246 606
rect 120 560 121 561
rect 122 560 123 561
rect 123 560 124 561
rect 125 560 126 561
rect 120 561 126 565
rect 120 565 121 566
rect 122 565 123 566
rect 123 565 124 566
rect 125 565 126 566
rect 800 480 801 481
rect 802 480 803 481
rect 803 480 804 481
rect 805 480 806 481
rect 800 481 806 485
rect 800 485 801 486
rect 802 485 803 486
rect 803 485 804 486
rect 805 485 806 486
rect 620 580 621 581
rect 622 580 623 581
rect 623 580 624 581
rect 625 580 626 581
rect 620 581 626 585
rect 620 585 621 586
rect 622 585 623 586
rect 623 585 624 586
rect 625 585 626 586
rect 780 560 781 561
rect 782 560 783 561
rect 783 560 784 561
rect 785 560 786 561
rect 780 561 786 565
rect 780 565 781 566
rect 782 565 783 566
rect 783 565 784 566
rect 785 565 786 566
rect 840 480 841 481
rect 842 480 843 481
rect 843 480 844 481
rect 845 480 846 481
rect 840 481 846 485
rect 840 485 841 486
rect 842 485 843 486
rect 843 485 844 486
rect 845 485 846 486
rect 600 480 601 481
rect 602 480 603 481
rect 603 480 604 481
rect 605 480 606 481
rect 600 481 606 485
rect 600 485 601 486
rect 602 485 603 486
rect 603 485 604 486
rect 605 485 606 486
rect 520 800 521 801
rect 522 800 523 801
rect 523 800 524 801
rect 525 800 526 801
rect 520 801 526 805
rect 520 805 521 806
rect 522 805 523 806
rect 523 805 524 806
rect 525 805 526 806
rect 480 200 481 201
rect 482 200 483 201
rect 483 200 484 201
rect 485 200 486 201
rect 480 201 486 205
rect 480 205 481 206
rect 482 205 483 206
rect 483 205 484 206
rect 485 205 486 206
rect 560 200 561 201
rect 562 200 563 201
rect 563 200 564 201
rect 565 200 566 201
rect 560 201 566 205
rect 560 205 561 206
rect 562 205 563 206
rect 563 205 564 206
rect 565 205 566 206
rect 720 400 721 401
rect 722 400 723 401
rect 723 400 724 401
rect 725 400 726 401
rect 720 401 726 405
rect 720 405 721 406
rect 722 405 723 406
rect 723 405 724 406
rect 725 405 726 406
rect 280 420 281 421
rect 282 420 283 421
rect 283 420 284 421
rect 285 420 286 421
rect 280 421 286 425
rect 280 425 281 426
rect 282 425 283 426
rect 283 425 284 426
rect 285 425 286 426
rect 820 420 821 421
rect 822 420 823 421
rect 823 420 824 421
rect 825 420 826 421
rect 820 421 826 425
rect 820 425 821 426
rect 822 425 823 426
rect 823 425 824 426
rect 825 425 826 426
rect 600 240 601 241
rect 602 240 603 241
rect 603 240 604 241
rect 605 240 606 241
rect 600 241 606 245
rect 600 245 601 246
rect 602 245 603 246
rect 603 245 604 246
rect 605 245 606 246
rect 620 340 621 341
rect 622 340 623 341
rect 623 340 624 341
rect 625 340 626 341
rect 620 341 626 345
rect 620 345 621 346
rect 622 345 623 346
rect 623 345 624 346
rect 625 345 626 346
rect 580 180 581 181
rect 582 180 583 181
rect 583 180 584 181
rect 585 180 586 181
rect 580 181 586 185
rect 580 185 581 186
rect 582 185 583 186
rect 583 185 584 186
rect 585 185 586 186
rect 720 620 721 621
rect 722 620 723 621
rect 723 620 724 621
rect 725 620 726 621
rect 720 621 726 625
rect 720 625 721 626
rect 722 625 723 626
rect 723 625 724 626
rect 725 625 726 626
rect 460 360 461 361
rect 462 360 463 361
rect 463 360 464 361
rect 465 360 466 361
rect 460 361 466 365
rect 460 365 461 366
rect 462 365 463 366
rect 463 365 464 366
rect 465 365 466 366
rect 460 380 461 381
rect 462 380 463 381
rect 463 380 464 381
rect 465 380 466 381
rect 460 381 466 385
rect 460 385 461 386
rect 462 385 463 386
rect 463 385 464 386
rect 465 385 466 386
rect 780 400 781 401
rect 782 400 783 401
rect 783 400 784 401
rect 785 400 786 401
rect 780 401 786 405
rect 780 405 781 406
rect 782 405 783 406
rect 783 405 784 406
rect 785 405 786 406
rect 600 580 601 581
rect 602 580 603 581
rect 603 580 604 581
rect 605 580 606 581
rect 600 581 606 585
rect 600 585 601 586
rect 602 585 603 586
rect 603 585 604 586
rect 605 585 606 586
rect 760 340 761 341
rect 762 340 763 341
rect 763 340 764 341
rect 765 340 766 341
rect 760 341 766 345
rect 760 345 761 346
rect 762 345 763 346
rect 763 345 764 346
rect 765 345 766 346
rect 620 600 621 601
rect 622 600 623 601
rect 623 600 624 601
rect 625 600 626 601
rect 620 601 626 605
rect 620 605 621 606
rect 622 605 623 606
rect 623 605 624 606
rect 625 605 626 606
rect 560 820 561 821
rect 562 820 563 821
rect 563 820 564 821
rect 565 820 566 821
rect 560 821 566 825
rect 560 825 561 826
rect 562 825 563 826
rect 563 825 564 826
rect 565 825 566 826
rect 480 680 481 681
rect 482 680 483 681
rect 483 680 484 681
rect 485 680 486 681
rect 480 681 486 685
rect 480 685 481 686
rect 482 685 483 686
rect 483 685 484 686
rect 485 685 486 686
rect 340 520 341 521
rect 342 520 343 521
rect 343 520 344 521
rect 345 520 346 521
rect 340 521 346 525
rect 340 525 341 526
rect 342 525 343 526
rect 343 525 344 526
rect 345 525 346 526
rect 180 440 181 441
rect 182 440 183 441
rect 183 440 184 441
rect 185 440 186 441
rect 180 441 186 445
rect 180 445 181 446
rect 182 445 183 446
rect 183 445 184 446
rect 185 445 186 446
rect 780 580 781 581
rect 782 580 783 581
rect 783 580 784 581
rect 785 580 786 581
rect 780 581 786 585
rect 780 585 781 586
rect 782 585 783 586
rect 783 585 784 586
rect 785 585 786 586
rect 640 680 641 681
rect 642 680 643 681
rect 643 680 644 681
rect 645 680 646 681
rect 640 681 646 685
rect 640 685 641 686
rect 642 685 643 686
rect 643 685 644 686
rect 645 685 646 686
rect 700 320 701 321
rect 702 320 703 321
rect 703 320 704 321
rect 705 320 706 321
rect 700 321 706 325
rect 700 325 701 326
rect 702 325 703 326
rect 703 325 704 326
rect 705 325 706 326
rect 340 420 341 421
rect 342 420 343 421
rect 343 420 344 421
rect 345 420 346 421
rect 340 421 346 425
rect 340 425 341 426
rect 342 425 343 426
rect 343 425 344 426
rect 345 425 346 426
rect 840 600 841 601
rect 842 600 843 601
rect 843 600 844 601
rect 845 600 846 601
rect 840 601 846 605
rect 840 605 841 606
rect 842 605 843 606
rect 843 605 844 606
rect 845 605 846 606
rect 300 640 301 641
rect 302 640 303 641
rect 303 640 304 641
rect 305 640 306 641
rect 300 641 306 645
rect 300 645 301 646
rect 302 645 303 646
rect 303 645 304 646
rect 305 645 306 646
rect 500 640 501 641
rect 502 640 503 641
rect 503 640 504 641
rect 505 640 506 641
rect 500 641 506 645
rect 500 645 501 646
rect 502 645 503 646
rect 503 645 504 646
rect 505 645 506 646
rect 440 520 441 521
rect 442 520 443 521
rect 443 520 444 521
rect 445 520 446 521
rect 440 521 446 525
rect 440 525 441 526
rect 442 525 443 526
rect 443 525 444 526
rect 445 525 446 526
rect 320 560 321 561
rect 322 560 323 561
rect 323 560 324 561
rect 325 560 326 561
rect 320 561 326 565
rect 320 565 321 566
rect 322 565 323 566
rect 323 565 324 566
rect 325 565 326 566
rect 480 380 481 381
rect 482 380 483 381
rect 483 380 484 381
rect 485 380 486 381
rect 480 381 486 385
rect 480 385 481 386
rect 482 385 483 386
rect 483 385 484 386
rect 485 385 486 386
rect 700 480 701 481
rect 702 480 703 481
rect 703 480 704 481
rect 705 480 706 481
rect 700 481 706 485
rect 700 485 701 486
rect 702 485 703 486
rect 703 485 704 486
rect 705 485 706 486
rect 380 440 381 441
rect 382 440 383 441
rect 383 440 384 441
rect 385 440 386 441
rect 380 441 386 445
rect 380 445 381 446
rect 382 445 383 446
rect 383 445 384 446
rect 385 445 386 446
rect 460 240 461 241
rect 462 240 463 241
rect 463 240 464 241
rect 465 240 466 241
rect 460 241 466 245
rect 460 245 461 246
rect 462 245 463 246
rect 463 245 464 246
rect 465 245 466 246
rect 400 360 401 361
rect 402 360 403 361
rect 403 360 404 361
rect 405 360 406 361
rect 400 361 406 365
rect 400 365 401 366
rect 402 365 403 366
rect 403 365 404 366
rect 405 365 406 366
rect 600 720 601 721
rect 602 720 603 721
rect 603 720 604 721
rect 605 720 606 721
rect 600 721 606 725
rect 600 725 601 726
rect 602 725 603 726
rect 603 725 604 726
rect 605 725 606 726
rect 460 700 461 701
rect 462 700 463 701
rect 463 700 464 701
rect 465 700 466 701
rect 460 701 466 705
rect 460 705 461 706
rect 462 705 463 706
rect 463 705 464 706
rect 465 705 466 706
rect 480 560 481 561
rect 482 560 483 561
rect 483 560 484 561
rect 485 560 486 561
rect 480 561 486 565
rect 480 565 481 566
rect 482 565 483 566
rect 483 565 484 566
rect 485 565 486 566
rect 660 760 661 761
rect 662 760 663 761
rect 663 760 664 761
rect 665 760 666 761
rect 660 761 666 765
rect 660 765 661 766
rect 662 765 663 766
rect 663 765 664 766
rect 665 765 666 766
rect 380 740 381 741
rect 382 740 383 741
rect 383 740 384 741
rect 385 740 386 741
rect 380 741 386 745
rect 380 745 381 746
rect 382 745 383 746
rect 383 745 384 746
rect 385 745 386 746
rect 680 760 681 761
rect 682 760 683 761
rect 683 760 684 761
rect 685 760 686 761
rect 680 761 686 765
rect 680 765 681 766
rect 682 765 683 766
rect 683 765 684 766
rect 685 765 686 766
rect 640 240 641 241
rect 642 240 643 241
rect 643 240 644 241
rect 645 240 646 241
rect 640 241 646 245
rect 640 245 641 246
rect 642 245 643 246
rect 643 245 644 246
rect 645 245 646 246
rect 740 500 741 501
rect 742 500 743 501
rect 743 500 744 501
rect 745 500 746 501
rect 740 501 746 505
rect 740 505 741 506
rect 742 505 743 506
rect 743 505 744 506
rect 745 505 746 506
rect 380 700 381 701
rect 382 700 383 701
rect 383 700 384 701
rect 385 700 386 701
rect 380 701 386 705
rect 380 705 381 706
rect 382 705 383 706
rect 383 705 384 706
rect 385 705 386 706
rect 380 580 381 581
rect 382 580 383 581
rect 383 580 384 581
rect 385 580 386 581
rect 380 581 386 585
rect 380 585 381 586
rect 382 585 383 586
rect 383 585 384 586
rect 385 585 386 586
rect 720 340 721 341
rect 722 340 723 341
rect 723 340 724 341
rect 725 340 726 341
rect 720 341 726 345
rect 720 345 721 346
rect 722 345 723 346
rect 723 345 724 346
rect 725 345 726 346
rect 400 180 401 181
rect 402 180 403 181
rect 403 180 404 181
rect 405 180 406 181
rect 400 181 406 185
rect 400 185 401 186
rect 402 185 403 186
rect 403 185 404 186
rect 405 185 406 186
rect 380 560 381 561
rect 382 560 383 561
rect 383 560 384 561
rect 385 560 386 561
rect 380 561 386 565
rect 380 565 381 566
rect 382 565 383 566
rect 383 565 384 566
rect 385 565 386 566
rect 520 320 521 321
rect 522 320 523 321
rect 523 320 524 321
rect 525 320 526 321
rect 520 321 526 325
rect 520 325 521 326
rect 522 325 523 326
rect 523 325 524 326
rect 525 325 526 326
rect 680 300 681 301
rect 682 300 683 301
rect 683 300 684 301
rect 685 300 686 301
rect 680 301 686 305
rect 680 305 681 306
rect 682 305 683 306
rect 683 305 684 306
rect 685 305 686 306
rect 660 260 661 261
rect 662 260 663 261
rect 663 260 664 261
rect 665 260 666 261
rect 660 261 666 265
rect 660 265 661 266
rect 662 265 663 266
rect 663 265 664 266
rect 665 265 666 266
rect 460 200 461 201
rect 462 200 463 201
rect 463 200 464 201
rect 465 200 466 201
rect 460 201 466 205
rect 460 205 461 206
rect 462 205 463 206
rect 463 205 464 206
rect 465 205 466 206
rect 220 620 221 621
rect 222 620 223 621
rect 223 620 224 621
rect 225 620 226 621
rect 220 621 226 625
rect 220 625 221 626
rect 222 625 223 626
rect 223 625 224 626
rect 225 625 226 626
rect 380 820 381 821
rect 382 820 383 821
rect 383 820 384 821
rect 385 820 386 821
rect 380 821 386 825
rect 380 825 381 826
rect 382 825 383 826
rect 383 825 384 826
rect 385 825 386 826
rect 620 640 621 641
rect 622 640 623 641
rect 623 640 624 641
rect 625 640 626 641
rect 620 641 626 645
rect 620 645 621 646
rect 622 645 623 646
rect 623 645 624 646
rect 625 645 626 646
rect 420 440 421 441
rect 422 440 423 441
rect 423 440 424 441
rect 425 440 426 441
rect 420 441 426 445
rect 420 445 421 446
rect 422 445 423 446
rect 423 445 424 446
rect 425 445 426 446
rect 320 520 321 521
rect 322 520 323 521
rect 323 520 324 521
rect 325 520 326 521
rect 320 521 326 525
rect 320 525 321 526
rect 322 525 323 526
rect 323 525 324 526
rect 325 525 326 526
rect 400 580 401 581
rect 402 580 403 581
rect 403 580 404 581
rect 405 580 406 581
rect 400 581 406 585
rect 400 585 401 586
rect 402 585 403 586
rect 403 585 404 586
rect 405 585 406 586
rect 380 800 381 801
rect 382 800 383 801
rect 383 800 384 801
rect 385 800 386 801
rect 380 801 386 805
rect 380 805 381 806
rect 382 805 383 806
rect 383 805 384 806
rect 385 805 386 806
rect 600 600 601 601
rect 602 600 603 601
rect 603 600 604 601
rect 605 600 606 601
rect 600 601 606 605
rect 600 605 601 606
rect 602 605 603 606
rect 603 605 604 606
rect 605 605 606 606
rect 540 740 541 741
rect 542 740 543 741
rect 543 740 544 741
rect 545 740 546 741
rect 540 741 546 745
rect 540 745 541 746
rect 542 745 543 746
rect 543 745 544 746
rect 545 745 546 746
rect 480 620 481 621
rect 482 620 483 621
rect 483 620 484 621
rect 485 620 486 621
rect 480 621 486 625
rect 480 625 481 626
rect 482 625 483 626
rect 483 625 484 626
rect 485 625 486 626
rect 800 520 801 521
rect 802 520 803 521
rect 803 520 804 521
rect 805 520 806 521
rect 800 521 806 525
rect 800 525 801 526
rect 802 525 803 526
rect 803 525 804 526
rect 805 525 806 526
rect 560 680 561 681
rect 562 680 563 681
rect 563 680 564 681
rect 565 680 566 681
rect 560 681 566 685
rect 560 685 561 686
rect 562 685 563 686
rect 563 685 564 686
rect 565 685 566 686
rect 580 620 581 621
rect 582 620 583 621
rect 583 620 584 621
rect 585 620 586 621
rect 580 621 586 625
rect 580 625 581 626
rect 582 625 583 626
rect 583 625 584 626
rect 585 625 586 626
rect 240 400 241 401
rect 242 400 243 401
rect 243 400 244 401
rect 245 400 246 401
rect 240 401 246 405
rect 240 405 241 406
rect 242 405 243 406
rect 243 405 244 406
rect 245 405 246 406
rect 600 360 601 361
rect 602 360 603 361
rect 603 360 604 361
rect 605 360 606 361
rect 600 361 606 365
rect 600 365 601 366
rect 602 365 603 366
rect 603 365 604 366
rect 605 365 606 366
rect 520 880 521 881
rect 522 880 523 881
rect 523 880 524 881
rect 525 880 526 881
rect 520 881 526 885
rect 520 885 521 886
rect 522 885 523 886
rect 523 885 524 886
rect 525 885 526 886
rect 540 380 541 381
rect 542 380 543 381
rect 543 380 544 381
rect 545 380 546 381
rect 540 381 546 385
rect 540 385 541 386
rect 542 385 543 386
rect 543 385 544 386
rect 545 385 546 386
rect 220 580 221 581
rect 222 580 223 581
rect 223 580 224 581
rect 225 580 226 581
rect 220 581 226 585
rect 220 585 221 586
rect 222 585 223 586
rect 223 585 224 586
rect 225 585 226 586
rect 680 740 681 741
rect 682 740 683 741
rect 683 740 684 741
rect 685 740 686 741
rect 680 741 686 745
rect 680 745 681 746
rect 682 745 683 746
rect 683 745 684 746
rect 685 745 686 746
rect 400 480 401 481
rect 402 480 403 481
rect 403 480 404 481
rect 405 480 406 481
rect 400 481 406 485
rect 400 485 401 486
rect 402 485 403 486
rect 403 485 404 486
rect 405 485 406 486
rect 760 620 761 621
rect 762 620 763 621
rect 763 620 764 621
rect 765 620 766 621
rect 760 621 766 625
rect 760 625 761 626
rect 762 625 763 626
rect 763 625 764 626
rect 765 625 766 626
rect 600 760 601 761
rect 602 760 603 761
rect 603 760 604 761
rect 605 760 606 761
rect 600 761 606 765
rect 600 765 601 766
rect 602 765 603 766
rect 603 765 604 766
rect 605 765 606 766
rect 600 660 601 661
rect 602 660 603 661
rect 603 660 604 661
rect 605 660 606 661
rect 600 661 606 665
rect 600 665 601 666
rect 602 665 603 666
rect 603 665 604 666
rect 605 665 606 666
rect 460 760 461 761
rect 462 760 463 761
rect 463 760 464 761
rect 465 760 466 761
rect 460 761 466 765
rect 460 765 461 766
rect 462 765 463 766
rect 463 765 464 766
rect 465 765 466 766
rect 600 320 601 321
rect 602 320 603 321
rect 603 320 604 321
rect 605 320 606 321
rect 600 321 606 325
rect 600 325 601 326
rect 602 325 603 326
rect 603 325 604 326
rect 605 325 606 326
rect 700 380 701 381
rect 702 380 703 381
rect 703 380 704 381
rect 705 380 706 381
rect 700 381 706 385
rect 700 385 701 386
rect 702 385 703 386
rect 703 385 704 386
rect 705 385 706 386
rect 700 720 701 721
rect 702 720 703 721
rect 703 720 704 721
rect 705 720 706 721
rect 700 721 706 725
rect 700 725 701 726
rect 702 725 703 726
rect 703 725 704 726
rect 705 725 706 726
rect 680 780 681 781
rect 682 780 683 781
rect 683 780 684 781
rect 685 780 686 781
rect 680 781 686 785
rect 680 785 681 786
rect 682 785 683 786
rect 683 785 684 786
rect 685 785 686 786
rect 540 720 541 721
rect 542 720 543 721
rect 543 720 544 721
rect 545 720 546 721
rect 540 721 546 725
rect 540 725 541 726
rect 542 725 543 726
rect 543 725 544 726
rect 545 725 546 726
rect 280 660 281 661
rect 282 660 283 661
rect 283 660 284 661
rect 285 660 286 661
rect 280 661 286 665
rect 280 665 281 666
rect 282 665 283 666
rect 283 665 284 666
rect 285 665 286 666
rect 760 440 761 441
rect 762 440 763 441
rect 763 440 764 441
rect 765 440 766 441
rect 760 441 766 445
rect 760 445 761 446
rect 762 445 763 446
rect 763 445 764 446
rect 765 445 766 446
rect 500 500 501 501
rect 502 500 503 501
rect 503 500 504 501
rect 505 500 506 501
rect 500 501 506 505
rect 500 505 501 506
rect 502 505 503 506
rect 503 505 504 506
rect 505 505 506 506
rect 240 460 241 461
rect 242 460 243 461
rect 243 460 244 461
rect 245 460 246 461
rect 240 461 246 465
rect 240 465 241 466
rect 242 465 243 466
rect 243 465 244 466
rect 245 465 246 466
rect 320 400 321 401
rect 322 400 323 401
rect 323 400 324 401
rect 325 400 326 401
rect 320 401 326 405
rect 320 405 321 406
rect 322 405 323 406
rect 323 405 324 406
rect 325 405 326 406
rect 540 860 541 861
rect 542 860 543 861
rect 543 860 544 861
rect 545 860 546 861
rect 540 861 546 865
rect 540 865 541 866
rect 542 865 543 866
rect 543 865 544 866
rect 545 865 546 866
rect 260 420 261 421
rect 262 420 263 421
rect 263 420 264 421
rect 265 420 266 421
rect 260 421 266 425
rect 260 425 261 426
rect 262 425 263 426
rect 263 425 264 426
rect 265 425 266 426
rect 680 620 681 621
rect 682 620 683 621
rect 683 620 684 621
rect 685 620 686 621
rect 680 621 686 625
rect 680 625 681 626
rect 682 625 683 626
rect 683 625 684 626
rect 685 625 686 626
rect 320 300 321 301
rect 322 300 323 301
rect 323 300 324 301
rect 325 300 326 301
rect 320 301 326 305
rect 320 305 321 306
rect 322 305 323 306
rect 323 305 324 306
rect 325 305 326 306
rect 640 660 641 661
rect 642 660 643 661
rect 643 660 644 661
rect 645 660 646 661
rect 640 661 646 665
rect 640 665 641 666
rect 642 665 643 666
rect 643 665 644 666
rect 645 665 646 666
rect 660 720 661 721
rect 662 720 663 721
rect 663 720 664 721
rect 665 720 666 721
rect 660 721 666 725
rect 660 725 661 726
rect 662 725 663 726
rect 663 725 664 726
rect 665 725 666 726
rect 580 500 581 501
rect 582 500 583 501
rect 583 500 584 501
rect 585 500 586 501
rect 580 501 586 505
rect 580 505 581 506
rect 582 505 583 506
rect 583 505 584 506
rect 585 505 586 506
rect 440 480 441 481
rect 442 480 443 481
rect 443 480 444 481
rect 445 480 446 481
rect 440 481 446 485
rect 440 485 441 486
rect 442 485 443 486
rect 443 485 444 486
rect 445 485 446 486
rect 680 800 681 801
rect 682 800 683 801
rect 683 800 684 801
rect 685 800 686 801
rect 680 801 686 805
rect 680 805 681 806
rect 682 805 683 806
rect 683 805 684 806
rect 685 805 686 806
rect 620 360 621 361
rect 622 360 623 361
rect 623 360 624 361
rect 625 360 626 361
rect 620 361 626 365
rect 620 365 621 366
rect 622 365 623 366
rect 623 365 624 366
rect 625 365 626 366
rect 500 480 501 481
rect 502 480 503 481
rect 503 480 504 481
rect 505 480 506 481
rect 500 481 506 485
rect 500 485 501 486
rect 502 485 503 486
rect 503 485 504 486
rect 505 485 506 486
rect 280 700 281 701
rect 282 700 283 701
rect 283 700 284 701
rect 285 700 286 701
rect 280 701 286 705
rect 280 705 281 706
rect 282 705 283 706
rect 283 705 284 706
rect 285 705 286 706
rect 200 600 201 601
rect 202 600 203 601
rect 203 600 204 601
rect 205 600 206 601
rect 200 601 206 605
rect 200 605 201 606
rect 202 605 203 606
rect 203 605 204 606
rect 205 605 206 606
rect 760 680 761 681
rect 762 680 763 681
rect 763 680 764 681
rect 765 680 766 681
rect 760 681 766 685
rect 760 685 761 686
rect 762 685 763 686
rect 763 685 764 686
rect 765 685 766 686
rect 580 540 581 541
rect 582 540 583 541
rect 583 540 584 541
rect 585 540 586 541
rect 580 541 586 545
rect 580 545 581 546
rect 582 545 583 546
rect 583 545 584 546
rect 585 545 586 546
rect 120 540 121 541
rect 122 540 123 541
rect 123 540 124 541
rect 125 540 126 541
rect 120 541 126 545
rect 120 545 121 546
rect 122 545 123 546
rect 123 545 124 546
rect 125 545 126 546
rect 180 600 181 601
rect 182 600 183 601
rect 183 600 184 601
rect 185 600 186 601
rect 180 601 186 605
rect 180 605 181 606
rect 182 605 183 606
rect 183 605 184 606
rect 185 605 186 606
rect 520 380 521 381
rect 522 380 523 381
rect 523 380 524 381
rect 525 380 526 381
rect 520 381 526 385
rect 520 385 521 386
rect 522 385 523 386
rect 523 385 524 386
rect 525 385 526 386
rect 500 440 501 441
rect 502 440 503 441
rect 503 440 504 441
rect 505 440 506 441
rect 500 441 506 445
rect 500 445 501 446
rect 502 445 503 446
rect 503 445 504 446
rect 505 445 506 446
rect 340 280 341 281
rect 342 280 343 281
rect 343 280 344 281
rect 345 280 346 281
rect 340 281 346 285
rect 340 285 341 286
rect 342 285 343 286
rect 343 285 344 286
rect 345 285 346 286
rect 440 420 441 421
rect 442 420 443 421
rect 443 420 444 421
rect 445 420 446 421
rect 440 421 446 425
rect 440 425 441 426
rect 442 425 443 426
rect 443 425 444 426
rect 445 425 446 426
rect 740 540 741 541
rect 742 540 743 541
rect 743 540 744 541
rect 745 540 746 541
rect 740 541 746 545
rect 740 545 741 546
rect 742 545 743 546
rect 743 545 744 546
rect 745 545 746 546
rect 540 880 541 881
rect 542 880 543 881
rect 543 880 544 881
rect 545 880 546 881
rect 540 881 546 885
rect 540 885 541 886
rect 542 885 543 886
rect 543 885 544 886
rect 545 885 546 886
rect 460 280 461 281
rect 462 280 463 281
rect 463 280 464 281
rect 465 280 466 281
rect 460 281 466 285
rect 460 285 461 286
rect 462 285 463 286
rect 463 285 464 286
rect 465 285 466 286
rect 380 540 381 541
rect 382 540 383 541
rect 383 540 384 541
rect 385 540 386 541
rect 380 541 386 545
rect 380 545 381 546
rect 382 545 383 546
rect 383 545 384 546
rect 385 545 386 546
rect 680 540 681 541
rect 682 540 683 541
rect 683 540 684 541
rect 685 540 686 541
rect 680 541 686 545
rect 680 545 681 546
rect 682 545 683 546
rect 683 545 684 546
rect 685 545 686 546
rect 500 300 501 301
rect 502 300 503 301
rect 503 300 504 301
rect 505 300 506 301
rect 500 301 506 305
rect 500 305 501 306
rect 502 305 503 306
rect 503 305 504 306
rect 505 305 506 306
rect 360 320 361 321
rect 362 320 363 321
rect 363 320 364 321
rect 365 320 366 321
rect 360 321 366 325
rect 360 325 361 326
rect 362 325 363 326
rect 363 325 364 326
rect 365 325 366 326
rect 520 340 521 341
rect 522 340 523 341
rect 523 340 524 341
rect 525 340 526 341
rect 520 341 526 345
rect 520 345 521 346
rect 522 345 523 346
rect 523 345 524 346
rect 525 345 526 346
rect 680 320 681 321
rect 682 320 683 321
rect 683 320 684 321
rect 685 320 686 321
rect 680 321 686 325
rect 680 325 681 326
rect 682 325 683 326
rect 683 325 684 326
rect 685 325 686 326
rect 540 700 541 701
rect 542 700 543 701
rect 543 700 544 701
rect 545 700 546 701
rect 540 701 546 705
rect 540 705 541 706
rect 542 705 543 706
rect 543 705 544 706
rect 545 705 546 706
rect 420 620 421 621
rect 422 620 423 621
rect 423 620 424 621
rect 425 620 426 621
rect 420 621 426 625
rect 420 625 421 626
rect 422 625 423 626
rect 423 625 424 626
rect 425 625 426 626
rect 660 560 661 561
rect 662 560 663 561
rect 663 560 664 561
rect 665 560 666 561
rect 660 561 666 565
rect 660 565 661 566
rect 662 565 663 566
rect 663 565 664 566
rect 665 565 666 566
rect 540 300 541 301
rect 542 300 543 301
rect 543 300 544 301
rect 545 300 546 301
rect 540 301 546 305
rect 540 305 541 306
rect 542 305 543 306
rect 543 305 544 306
rect 545 305 546 306
rect 540 800 541 801
rect 542 800 543 801
rect 543 800 544 801
rect 545 800 546 801
rect 540 801 546 805
rect 540 805 541 806
rect 542 805 543 806
rect 543 805 544 806
rect 545 805 546 806
rect 300 460 301 461
rect 302 460 303 461
rect 303 460 304 461
rect 305 460 306 461
rect 300 461 306 465
rect 300 465 301 466
rect 302 465 303 466
rect 303 465 304 466
rect 305 465 306 466
rect 580 600 581 601
rect 582 600 583 601
rect 583 600 584 601
rect 585 600 586 601
rect 580 601 586 605
rect 580 605 581 606
rect 582 605 583 606
rect 583 605 584 606
rect 585 605 586 606
rect 380 780 381 781
rect 382 780 383 781
rect 383 780 384 781
rect 385 780 386 781
rect 380 781 386 785
rect 380 785 381 786
rect 382 785 383 786
rect 383 785 384 786
rect 385 785 386 786
rect 480 480 481 481
rect 482 480 483 481
rect 483 480 484 481
rect 485 480 486 481
rect 480 481 486 485
rect 480 485 481 486
rect 482 485 483 486
rect 483 485 484 486
rect 485 485 486 486
rect 400 400 401 401
rect 402 400 403 401
rect 403 400 404 401
rect 405 400 406 401
rect 400 401 406 405
rect 400 405 401 406
rect 402 405 403 406
rect 403 405 404 406
rect 405 405 406 406
rect 580 300 581 301
rect 582 300 583 301
rect 583 300 584 301
rect 585 300 586 301
rect 580 301 586 305
rect 580 305 581 306
rect 582 305 583 306
rect 583 305 584 306
rect 585 305 586 306
rect 660 420 661 421
rect 662 420 663 421
rect 663 420 664 421
rect 665 420 666 421
rect 660 421 666 425
rect 660 425 661 426
rect 662 425 663 426
rect 663 425 664 426
rect 665 425 666 426
rect 200 400 201 401
rect 202 400 203 401
rect 203 400 204 401
rect 205 400 206 401
rect 200 401 206 405
rect 200 405 201 406
rect 202 405 203 406
rect 203 405 204 406
rect 205 405 206 406
rect 520 240 521 241
rect 522 240 523 241
rect 523 240 524 241
rect 525 240 526 241
rect 520 241 526 245
rect 520 245 521 246
rect 522 245 523 246
rect 523 245 524 246
rect 525 245 526 246
rect 340 660 341 661
rect 342 660 343 661
rect 343 660 344 661
rect 345 660 346 661
rect 340 661 346 665
rect 340 665 341 666
rect 342 665 343 666
rect 343 665 344 666
rect 345 665 346 666
rect 800 660 801 661
rect 802 660 803 661
rect 803 660 804 661
rect 805 660 806 661
rect 800 661 806 665
rect 800 665 801 666
rect 802 665 803 666
rect 803 665 804 666
rect 805 665 806 666
rect 300 520 301 521
rect 302 520 303 521
rect 303 520 304 521
rect 305 520 306 521
rect 300 521 306 525
rect 300 525 301 526
rect 302 525 303 526
rect 303 525 304 526
rect 305 525 306 526
rect 660 300 661 301
rect 662 300 663 301
rect 663 300 664 301
rect 665 300 666 301
rect 660 301 666 305
rect 660 305 661 306
rect 662 305 663 306
rect 663 305 664 306
rect 665 305 666 306
rect 600 500 601 501
rect 602 500 603 501
rect 603 500 604 501
rect 605 500 606 501
rect 600 501 606 505
rect 600 505 601 506
rect 602 505 603 506
rect 603 505 604 506
rect 605 505 606 506
rect 340 240 341 241
rect 342 240 343 241
rect 343 240 344 241
rect 345 240 346 241
rect 340 241 346 245
rect 340 245 341 246
rect 342 245 343 246
rect 343 245 344 246
rect 345 245 346 246
rect 740 420 741 421
rect 742 420 743 421
rect 743 420 744 421
rect 745 420 746 421
rect 740 421 746 425
rect 740 425 741 426
rect 742 425 743 426
rect 743 425 744 426
rect 745 425 746 426
rect 580 860 581 861
rect 582 860 583 861
rect 583 860 584 861
rect 585 860 586 861
rect 580 861 586 865
rect 580 865 581 866
rect 582 865 583 866
rect 583 865 584 866
rect 585 865 586 866
rect 200 460 201 461
rect 202 460 203 461
rect 203 460 204 461
rect 205 460 206 461
rect 200 461 206 465
rect 200 465 201 466
rect 202 465 203 466
rect 203 465 204 466
rect 205 465 206 466
rect 720 380 721 381
rect 722 380 723 381
rect 723 380 724 381
rect 725 380 726 381
rect 720 381 726 385
rect 720 385 721 386
rect 722 385 723 386
rect 723 385 724 386
rect 725 385 726 386
rect 420 760 421 761
rect 422 760 423 761
rect 423 760 424 761
rect 425 760 426 761
rect 420 761 426 765
rect 420 765 421 766
rect 422 765 423 766
rect 423 765 424 766
rect 425 765 426 766
rect 640 760 641 761
rect 642 760 643 761
rect 643 760 644 761
rect 645 760 646 761
rect 640 761 646 765
rect 640 765 641 766
rect 642 765 643 766
rect 643 765 644 766
rect 645 765 646 766
rect 580 380 581 381
rect 582 380 583 381
rect 583 380 584 381
rect 585 380 586 381
rect 580 381 586 385
rect 580 385 581 386
rect 582 385 583 386
rect 583 385 584 386
rect 585 385 586 386
rect 560 840 561 841
rect 562 840 563 841
rect 563 840 564 841
rect 565 840 566 841
rect 560 841 566 845
rect 560 845 561 846
rect 562 845 563 846
rect 563 845 564 846
rect 565 845 566 846
rect 380 620 381 621
rect 382 620 383 621
rect 383 620 384 621
rect 385 620 386 621
rect 380 621 386 625
rect 380 625 381 626
rect 382 625 383 626
rect 383 625 384 626
rect 385 625 386 626
rect 680 460 681 461
rect 682 460 683 461
rect 683 460 684 461
rect 685 460 686 461
rect 680 461 686 465
rect 680 465 681 466
rect 682 465 683 466
rect 683 465 684 466
rect 685 465 686 466
rect 460 560 461 561
rect 462 560 463 561
rect 463 560 464 561
rect 465 560 466 561
rect 460 561 466 565
rect 460 565 461 566
rect 462 565 463 566
rect 463 565 464 566
rect 465 565 466 566
rect 620 320 621 321
rect 622 320 623 321
rect 623 320 624 321
rect 625 320 626 321
rect 620 321 626 325
rect 620 325 621 326
rect 622 325 623 326
rect 623 325 624 326
rect 625 325 626 326
rect 500 360 501 361
rect 502 360 503 361
rect 503 360 504 361
rect 505 360 506 361
rect 500 361 506 365
rect 500 365 501 366
rect 502 365 503 366
rect 503 365 504 366
rect 505 365 506 366
rect 600 300 601 301
rect 602 300 603 301
rect 603 300 604 301
rect 605 300 606 301
rect 600 301 606 305
rect 600 305 601 306
rect 602 305 603 306
rect 603 305 604 306
rect 605 305 606 306
rect 440 400 441 401
rect 442 400 443 401
rect 443 400 444 401
rect 445 400 446 401
rect 440 401 446 405
rect 440 405 441 406
rect 442 405 443 406
rect 443 405 444 406
rect 445 405 446 406
rect 400 720 401 721
rect 402 720 403 721
rect 403 720 404 721
rect 405 720 406 721
rect 400 721 406 725
rect 400 725 401 726
rect 402 725 403 726
rect 403 725 404 726
rect 405 725 406 726
rect 880 580 881 581
rect 882 580 883 581
rect 883 580 884 581
rect 885 580 886 581
rect 880 581 886 585
rect 880 585 881 586
rect 882 585 883 586
rect 883 585 884 586
rect 885 585 886 586
rect 320 740 321 741
rect 322 740 323 741
rect 323 740 324 741
rect 325 740 326 741
rect 320 741 326 745
rect 320 745 321 746
rect 322 745 323 746
rect 323 745 324 746
rect 325 745 326 746
rect 580 840 581 841
rect 582 840 583 841
rect 583 840 584 841
rect 585 840 586 841
rect 580 841 586 845
rect 580 845 581 846
rect 582 845 583 846
rect 583 845 584 846
rect 585 845 586 846
rect 520 480 521 481
rect 522 480 523 481
rect 523 480 524 481
rect 525 480 526 481
rect 520 481 526 485
rect 520 485 521 486
rect 522 485 523 486
rect 523 485 524 486
rect 525 485 526 486
rect 300 760 301 761
rect 302 760 303 761
rect 303 760 304 761
rect 305 760 306 761
rect 300 761 306 765
rect 300 765 301 766
rect 302 765 303 766
rect 303 765 304 766
rect 305 765 306 766
rect 840 520 841 521
rect 842 520 843 521
rect 843 520 844 521
rect 845 520 846 521
rect 840 521 846 525
rect 840 525 841 526
rect 842 525 843 526
rect 843 525 844 526
rect 845 525 846 526
rect 400 200 401 201
rect 402 200 403 201
rect 403 200 404 201
rect 405 200 406 201
rect 400 201 406 205
rect 400 205 401 206
rect 402 205 403 206
rect 403 205 404 206
rect 405 205 406 206
rect 560 380 561 381
rect 562 380 563 381
rect 563 380 564 381
rect 565 380 566 381
rect 560 381 566 385
rect 560 385 561 386
rect 562 385 563 386
rect 563 385 564 386
rect 565 385 566 386
rect 360 240 361 241
rect 362 240 363 241
rect 363 240 364 241
rect 365 240 366 241
rect 360 241 366 245
rect 360 245 361 246
rect 362 245 363 246
rect 363 245 364 246
rect 365 245 366 246
rect 380 500 381 501
rect 382 500 383 501
rect 383 500 384 501
rect 385 500 386 501
rect 380 501 386 505
rect 380 505 381 506
rect 382 505 383 506
rect 383 505 384 506
rect 385 505 386 506
rect 560 520 561 521
rect 562 520 563 521
rect 563 520 564 521
rect 565 520 566 521
rect 560 521 566 525
rect 560 525 561 526
rect 562 525 563 526
rect 563 525 564 526
rect 565 525 566 526
rect 160 640 161 641
rect 162 640 163 641
rect 163 640 164 641
rect 165 640 166 641
rect 160 641 166 645
rect 160 645 161 646
rect 162 645 163 646
rect 163 645 164 646
rect 165 645 166 646
rect 580 460 581 461
rect 582 460 583 461
rect 583 460 584 461
rect 585 460 586 461
rect 580 461 586 465
rect 580 465 581 466
rect 582 465 583 466
rect 583 465 584 466
rect 585 465 586 466
rect 480 500 481 501
rect 482 500 483 501
rect 483 500 484 501
rect 485 500 486 501
rect 480 501 486 505
rect 480 505 481 506
rect 482 505 483 506
rect 483 505 484 506
rect 485 505 486 506
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect 660 680 661 681
rect 662 680 663 681
rect 663 680 664 681
rect 665 680 666 681
rect 660 681 666 685
rect 660 685 661 686
rect 662 685 663 686
rect 663 685 664 686
rect 665 685 666 686
rect 480 600 481 601
rect 482 600 483 601
rect 483 600 484 601
rect 485 600 486 601
rect 480 601 486 605
rect 480 605 481 606
rect 482 605 483 606
rect 483 605 484 606
rect 485 605 486 606
rect 240 720 241 721
rect 242 720 243 721
rect 243 720 244 721
rect 245 720 246 721
rect 240 721 246 725
rect 240 725 241 726
rect 242 725 243 726
rect 243 725 244 726
rect 245 725 246 726
rect 340 360 341 361
rect 342 360 343 361
rect 343 360 344 361
rect 345 360 346 361
rect 340 361 346 365
rect 340 365 341 366
rect 342 365 343 366
rect 343 365 344 366
rect 345 365 346 366
rect 360 640 361 641
rect 362 640 363 641
rect 363 640 364 641
rect 365 640 366 641
rect 360 641 366 645
rect 360 645 361 646
rect 362 645 363 646
rect 363 645 364 646
rect 365 645 366 646
rect 400 680 401 681
rect 402 680 403 681
rect 403 680 404 681
rect 405 680 406 681
rect 400 681 406 685
rect 400 685 401 686
rect 402 685 403 686
rect 403 685 404 686
rect 405 685 406 686
rect 580 360 581 361
rect 582 360 583 361
rect 583 360 584 361
rect 585 360 586 361
rect 580 361 586 365
rect 580 365 581 366
rect 582 365 583 366
rect 583 365 584 366
rect 585 365 586 366
rect 620 280 621 281
rect 622 280 623 281
rect 623 280 624 281
rect 625 280 626 281
rect 620 281 626 285
rect 620 285 621 286
rect 622 285 623 286
rect 623 285 624 286
rect 625 285 626 286
rect 600 180 601 181
rect 602 180 603 181
rect 603 180 604 181
rect 605 180 606 181
rect 600 181 606 185
rect 600 185 601 186
rect 602 185 603 186
rect 603 185 604 186
rect 605 185 606 186
rect 680 640 681 641
rect 682 640 683 641
rect 683 640 684 641
rect 685 640 686 641
rect 680 641 686 645
rect 680 645 681 646
rect 682 645 683 646
rect 683 645 684 646
rect 685 645 686 646
rect 500 160 501 161
rect 502 160 503 161
rect 503 160 504 161
rect 505 160 506 161
rect 500 161 506 165
rect 500 165 501 166
rect 502 165 503 166
rect 503 165 504 166
rect 505 165 506 166
rect 560 340 561 341
rect 562 340 563 341
rect 563 340 564 341
rect 565 340 566 341
rect 560 341 566 345
rect 560 345 561 346
rect 562 345 563 346
rect 563 345 564 346
rect 565 345 566 346
rect 680 340 681 341
rect 682 340 683 341
rect 683 340 684 341
rect 685 340 686 341
rect 680 341 686 345
rect 680 345 681 346
rect 682 345 683 346
rect 683 345 684 346
rect 685 345 686 346
rect 520 900 521 901
rect 522 900 523 901
rect 523 900 524 901
rect 525 900 526 901
rect 520 901 526 905
rect 520 905 521 906
rect 522 905 523 906
rect 523 905 524 906
rect 525 905 526 906
rect 580 280 581 281
rect 582 280 583 281
rect 583 280 584 281
rect 585 280 586 281
rect 580 281 586 285
rect 580 285 581 286
rect 582 285 583 286
rect 583 285 584 286
rect 585 285 586 286
rect 560 780 561 781
rect 562 780 563 781
rect 563 780 564 781
rect 565 780 566 781
rect 560 781 566 785
rect 560 785 561 786
rect 562 785 563 786
rect 563 785 564 786
rect 565 785 566 786
rect 400 380 401 381
rect 402 380 403 381
rect 403 380 404 381
rect 405 380 406 381
rect 400 381 406 385
rect 400 385 401 386
rect 402 385 403 386
rect 403 385 404 386
rect 405 385 406 386
rect 280 360 281 361
rect 282 360 283 361
rect 283 360 284 361
rect 285 360 286 361
rect 280 361 286 365
rect 280 365 281 366
rect 282 365 283 366
rect 283 365 284 366
rect 285 365 286 366
rect 440 640 441 641
rect 442 640 443 641
rect 443 640 444 641
rect 445 640 446 641
rect 440 641 446 645
rect 440 645 441 646
rect 442 645 443 646
rect 443 645 444 646
rect 445 645 446 646
rect 560 180 561 181
rect 562 180 563 181
rect 563 180 564 181
rect 565 180 566 181
rect 560 181 566 185
rect 560 185 561 186
rect 562 185 563 186
rect 563 185 564 186
rect 565 185 566 186
rect 780 460 781 461
rect 782 460 783 461
rect 783 460 784 461
rect 785 460 786 461
rect 780 461 786 465
rect 780 465 781 466
rect 782 465 783 466
rect 783 465 784 466
rect 785 465 786 466
rect 860 440 861 441
rect 862 440 863 441
rect 863 440 864 441
rect 865 440 866 441
rect 860 441 866 445
rect 860 445 861 446
rect 862 445 863 446
rect 863 445 864 446
rect 865 445 866 446
rect 780 600 781 601
rect 782 600 783 601
rect 783 600 784 601
rect 785 600 786 601
rect 780 601 786 605
rect 780 605 781 606
rect 782 605 783 606
rect 783 605 784 606
rect 785 605 786 606
rect 360 460 361 461
rect 362 460 363 461
rect 363 460 364 461
rect 365 460 366 461
rect 360 461 366 465
rect 360 465 361 466
rect 362 465 363 466
rect 363 465 364 466
rect 365 465 366 466
rect 400 520 401 521
rect 402 520 403 521
rect 403 520 404 521
rect 405 520 406 521
rect 400 521 406 525
rect 400 525 401 526
rect 402 525 403 526
rect 403 525 404 526
rect 405 525 406 526
rect 740 340 741 341
rect 742 340 743 341
rect 743 340 744 341
rect 745 340 746 341
rect 740 341 746 345
rect 740 345 741 346
rect 742 345 743 346
rect 743 345 744 346
rect 745 345 746 346
rect 820 540 821 541
rect 822 540 823 541
rect 823 540 824 541
rect 825 540 826 541
rect 820 541 826 545
rect 820 545 821 546
rect 822 545 823 546
rect 823 545 824 546
rect 825 545 826 546
rect 440 260 441 261
rect 442 260 443 261
rect 443 260 444 261
rect 445 260 446 261
rect 440 261 446 265
rect 440 265 441 266
rect 442 265 443 266
rect 443 265 444 266
rect 445 265 446 266
rect 340 460 341 461
rect 342 460 343 461
rect 343 460 344 461
rect 345 460 346 461
rect 340 461 346 465
rect 340 465 341 466
rect 342 465 343 466
rect 343 465 344 466
rect 345 465 346 466
rect 660 400 661 401
rect 662 400 663 401
rect 663 400 664 401
rect 665 400 666 401
rect 660 401 666 405
rect 660 405 661 406
rect 662 405 663 406
rect 663 405 664 406
rect 665 405 666 406
rect 560 560 561 561
rect 562 560 563 561
rect 563 560 564 561
rect 565 560 566 561
rect 560 561 566 565
rect 560 565 561 566
rect 562 565 563 566
rect 563 565 564 566
rect 565 565 566 566
rect 600 260 601 261
rect 602 260 603 261
rect 603 260 604 261
rect 605 260 606 261
rect 600 261 606 265
rect 600 265 601 266
rect 602 265 603 266
rect 603 265 604 266
rect 605 265 606 266
rect 780 480 781 481
rect 782 480 783 481
rect 783 480 784 481
rect 785 480 786 481
rect 780 481 786 485
rect 780 485 781 486
rect 782 485 783 486
rect 783 485 784 486
rect 785 485 786 486
rect 440 220 441 221
rect 442 220 443 221
rect 443 220 444 221
rect 445 220 446 221
rect 440 221 446 225
rect 440 225 441 226
rect 442 225 443 226
rect 443 225 444 226
rect 445 225 446 226
rect 200 560 201 561
rect 202 560 203 561
rect 203 560 204 561
rect 205 560 206 561
rect 200 561 206 565
rect 200 565 201 566
rect 202 565 203 566
rect 203 565 204 566
rect 205 565 206 566
rect 180 460 181 461
rect 182 460 183 461
rect 183 460 184 461
rect 185 460 186 461
rect 180 461 186 465
rect 180 465 181 466
rect 182 465 183 466
rect 183 465 184 466
rect 185 465 186 466
rect 300 780 301 781
rect 302 780 303 781
rect 303 780 304 781
rect 305 780 306 781
rect 300 781 306 785
rect 300 785 301 786
rect 302 785 303 786
rect 303 785 304 786
rect 305 785 306 786
rect 660 700 661 701
rect 662 700 663 701
rect 663 700 664 701
rect 665 700 666 701
rect 660 701 666 705
rect 660 705 661 706
rect 662 705 663 706
rect 663 705 664 706
rect 665 705 666 706
rect 600 380 601 381
rect 602 380 603 381
rect 603 380 604 381
rect 605 380 606 381
rect 600 381 606 385
rect 600 385 601 386
rect 602 385 603 386
rect 603 385 604 386
rect 605 385 606 386
rect 620 240 621 241
rect 622 240 623 241
rect 623 240 624 241
rect 625 240 626 241
rect 620 241 626 245
rect 620 245 621 246
rect 622 245 623 246
rect 623 245 624 246
rect 625 245 626 246
rect 720 700 721 701
rect 722 700 723 701
rect 723 700 724 701
rect 725 700 726 701
rect 720 701 726 705
rect 720 705 721 706
rect 722 705 723 706
rect 723 705 724 706
rect 725 705 726 706
rect 420 300 421 301
rect 422 300 423 301
rect 423 300 424 301
rect 425 300 426 301
rect 420 301 426 305
rect 420 305 421 306
rect 422 305 423 306
rect 423 305 424 306
rect 425 305 426 306
rect 180 400 181 401
rect 182 400 183 401
rect 183 400 184 401
rect 185 400 186 401
rect 180 401 186 405
rect 180 405 181 406
rect 182 405 183 406
rect 183 405 184 406
rect 185 405 186 406
rect 420 240 421 241
rect 422 240 423 241
rect 423 240 424 241
rect 425 240 426 241
rect 420 241 426 245
rect 420 245 421 246
rect 422 245 423 246
rect 423 245 424 246
rect 425 245 426 246
rect 520 500 521 501
rect 522 500 523 501
rect 523 500 524 501
rect 525 500 526 501
rect 520 501 526 505
rect 520 505 521 506
rect 522 505 523 506
rect 523 505 524 506
rect 525 505 526 506
rect 680 420 681 421
rect 682 420 683 421
rect 683 420 684 421
rect 685 420 686 421
rect 680 421 686 425
rect 680 425 681 426
rect 682 425 683 426
rect 683 425 684 426
rect 685 425 686 426
rect 360 480 361 481
rect 362 480 363 481
rect 363 480 364 481
rect 365 480 366 481
rect 360 481 366 485
rect 360 485 361 486
rect 362 485 363 486
rect 363 485 364 486
rect 365 485 366 486
rect 760 580 761 581
rect 762 580 763 581
rect 763 580 764 581
rect 765 580 766 581
rect 760 581 766 585
rect 760 585 761 586
rect 762 585 763 586
rect 763 585 764 586
rect 765 585 766 586
rect 600 640 601 641
rect 602 640 603 641
rect 603 640 604 641
rect 605 640 606 641
rect 600 641 606 645
rect 600 645 601 646
rect 602 645 603 646
rect 603 645 604 646
rect 605 645 606 646
rect 300 400 301 401
rect 302 400 303 401
rect 303 400 304 401
rect 305 400 306 401
rect 300 401 306 405
rect 300 405 301 406
rect 302 405 303 406
rect 303 405 304 406
rect 305 405 306 406
rect 200 480 201 481
rect 202 480 203 481
rect 203 480 204 481
rect 205 480 206 481
rect 200 481 206 485
rect 200 485 201 486
rect 202 485 203 486
rect 203 485 204 486
rect 205 485 206 486
rect 660 480 661 481
rect 662 480 663 481
rect 663 480 664 481
rect 665 480 666 481
rect 660 481 666 485
rect 660 485 661 486
rect 662 485 663 486
rect 663 485 664 486
rect 665 485 666 486
rect 740 560 741 561
rect 742 560 743 561
rect 743 560 744 561
rect 745 560 746 561
rect 740 561 746 565
rect 740 565 741 566
rect 742 565 743 566
rect 743 565 744 566
rect 745 565 746 566
rect 720 600 721 601
rect 722 600 723 601
rect 723 600 724 601
rect 725 600 726 601
rect 720 601 726 605
rect 720 605 721 606
rect 722 605 723 606
rect 723 605 724 606
rect 725 605 726 606
rect 640 740 641 741
rect 642 740 643 741
rect 643 740 644 741
rect 645 740 646 741
rect 640 741 646 745
rect 640 745 641 746
rect 642 745 643 746
rect 643 745 644 746
rect 645 745 646 746
rect 300 340 301 341
rect 302 340 303 341
rect 303 340 304 341
rect 305 340 306 341
rect 300 341 306 345
rect 300 345 301 346
rect 302 345 303 346
rect 303 345 304 346
rect 305 345 306 346
rect 720 320 721 321
rect 722 320 723 321
rect 723 320 724 321
rect 725 320 726 321
rect 720 321 726 325
rect 720 325 721 326
rect 722 325 723 326
rect 723 325 724 326
rect 725 325 726 326
rect 240 740 241 741
rect 242 740 243 741
rect 243 740 244 741
rect 245 740 246 741
rect 240 741 246 745
rect 240 745 241 746
rect 242 745 243 746
rect 243 745 244 746
rect 245 745 246 746
rect 480 880 481 881
rect 482 880 483 881
rect 483 880 484 881
rect 485 880 486 881
rect 480 881 486 885
rect 480 885 481 886
rect 482 885 483 886
rect 483 885 484 886
rect 485 885 486 886
rect 560 440 561 441
rect 562 440 563 441
rect 563 440 564 441
rect 565 440 566 441
rect 560 441 566 445
rect 560 445 561 446
rect 562 445 563 446
rect 563 445 564 446
rect 565 445 566 446
rect 480 360 481 361
rect 482 360 483 361
rect 483 360 484 361
rect 485 360 486 361
rect 480 361 486 365
rect 480 365 481 366
rect 482 365 483 366
rect 483 365 484 366
rect 485 365 486 366
rect 600 540 601 541
rect 602 540 603 541
rect 603 540 604 541
rect 605 540 606 541
rect 600 541 606 545
rect 600 545 601 546
rect 602 545 603 546
rect 603 545 604 546
rect 605 545 606 546
rect 660 520 661 521
rect 662 520 663 521
rect 663 520 664 521
rect 665 520 666 521
rect 660 521 666 525
rect 660 525 661 526
rect 662 525 663 526
rect 663 525 664 526
rect 665 525 666 526
rect 360 360 361 361
rect 362 360 363 361
rect 363 360 364 361
rect 365 360 366 361
rect 360 361 366 365
rect 360 365 361 366
rect 362 365 363 366
rect 363 365 364 366
rect 365 365 366 366
rect 220 380 221 381
rect 222 380 223 381
rect 223 380 224 381
rect 225 380 226 381
rect 220 381 226 385
rect 220 385 221 386
rect 222 385 223 386
rect 223 385 224 386
rect 225 385 226 386
rect 820 620 821 621
rect 822 620 823 621
rect 823 620 824 621
rect 825 620 826 621
rect 820 621 826 625
rect 820 625 821 626
rect 822 625 823 626
rect 823 625 824 626
rect 825 625 826 626
rect 680 280 681 281
rect 682 280 683 281
rect 683 280 684 281
rect 685 280 686 281
rect 680 281 686 285
rect 680 285 681 286
rect 682 285 683 286
rect 683 285 684 286
rect 685 285 686 286
rect 360 680 361 681
rect 362 680 363 681
rect 363 680 364 681
rect 365 680 366 681
rect 360 681 366 685
rect 360 685 361 686
rect 362 685 363 686
rect 363 685 364 686
rect 365 685 366 686
rect 360 660 361 661
rect 362 660 363 661
rect 363 660 364 661
rect 365 660 366 661
rect 360 661 366 665
rect 360 665 361 666
rect 362 665 363 666
rect 363 665 364 666
rect 365 665 366 666
rect 160 460 161 461
rect 162 460 163 461
rect 163 460 164 461
rect 165 460 166 461
rect 160 461 166 465
rect 160 465 161 466
rect 162 465 163 466
rect 163 465 164 466
rect 165 465 166 466
rect 480 520 481 521
rect 482 520 483 521
rect 483 520 484 521
rect 485 520 486 521
rect 480 521 486 525
rect 480 525 481 526
rect 482 525 483 526
rect 483 525 484 526
rect 485 525 486 526
rect 360 500 361 501
rect 362 500 363 501
rect 363 500 364 501
rect 365 500 366 501
rect 360 501 366 505
rect 360 505 361 506
rect 362 505 363 506
rect 363 505 364 506
rect 365 505 366 506
rect 540 780 541 781
rect 542 780 543 781
rect 543 780 544 781
rect 545 780 546 781
rect 540 781 546 785
rect 540 785 541 786
rect 542 785 543 786
rect 543 785 544 786
rect 545 785 546 786
rect 560 120 561 121
rect 562 120 563 121
rect 563 120 564 121
rect 565 120 566 121
rect 560 121 566 125
rect 560 125 561 126
rect 562 125 563 126
rect 563 125 564 126
rect 565 125 566 126
rect 740 620 741 621
rect 742 620 743 621
rect 743 620 744 621
rect 745 620 746 621
rect 740 621 746 625
rect 740 625 741 626
rect 742 625 743 626
rect 743 625 744 626
rect 745 625 746 626
rect 540 360 541 361
rect 542 360 543 361
rect 543 360 544 361
rect 545 360 546 361
rect 540 361 546 365
rect 540 365 541 366
rect 542 365 543 366
rect 543 365 544 366
rect 545 365 546 366
rect 320 440 321 441
rect 322 440 323 441
rect 323 440 324 441
rect 325 440 326 441
rect 320 441 326 445
rect 320 445 321 446
rect 322 445 323 446
rect 323 445 324 446
rect 325 445 326 446
rect 660 460 661 461
rect 662 460 663 461
rect 663 460 664 461
rect 665 460 666 461
rect 660 461 666 465
rect 660 465 661 466
rect 662 465 663 466
rect 663 465 664 466
rect 665 465 666 466
rect 580 240 581 241
rect 582 240 583 241
rect 583 240 584 241
rect 585 240 586 241
rect 580 241 586 245
rect 580 245 581 246
rect 582 245 583 246
rect 583 245 584 246
rect 585 245 586 246
rect 460 820 461 821
rect 462 820 463 821
rect 463 820 464 821
rect 465 820 466 821
rect 460 821 466 825
rect 460 825 461 826
rect 462 825 463 826
rect 463 825 464 826
rect 465 825 466 826
rect 620 740 621 741
rect 622 740 623 741
rect 623 740 624 741
rect 625 740 626 741
rect 620 741 626 745
rect 620 745 621 746
rect 622 745 623 746
rect 623 745 624 746
rect 625 745 626 746
rect 660 660 661 661
rect 662 660 663 661
rect 663 660 664 661
rect 665 660 666 661
rect 660 661 666 665
rect 660 665 661 666
rect 662 665 663 666
rect 663 665 664 666
rect 665 665 666 666
rect 500 320 501 321
rect 502 320 503 321
rect 503 320 504 321
rect 505 320 506 321
rect 500 321 506 325
rect 500 325 501 326
rect 502 325 503 326
rect 503 325 504 326
rect 505 325 506 326
rect 700 460 701 461
rect 702 460 703 461
rect 703 460 704 461
rect 705 460 706 461
rect 700 461 706 465
rect 700 465 701 466
rect 702 465 703 466
rect 703 465 704 466
rect 705 465 706 466
rect 660 600 661 601
rect 662 600 663 601
rect 663 600 664 601
rect 665 600 666 601
rect 660 601 666 605
rect 660 605 661 606
rect 662 605 663 606
rect 663 605 664 606
rect 665 605 666 606
rect 440 700 441 701
rect 442 700 443 701
rect 443 700 444 701
rect 445 700 446 701
rect 440 701 446 705
rect 440 705 441 706
rect 442 705 443 706
rect 443 705 444 706
rect 445 705 446 706
rect 240 320 241 321
rect 242 320 243 321
rect 243 320 244 321
rect 245 320 246 321
rect 240 321 246 325
rect 240 325 241 326
rect 242 325 243 326
rect 243 325 244 326
rect 245 325 246 326
rect 320 660 321 661
rect 322 660 323 661
rect 323 660 324 661
rect 325 660 326 661
rect 320 661 326 665
rect 320 665 321 666
rect 322 665 323 666
rect 323 665 324 666
rect 325 665 326 666
rect 360 720 361 721
rect 362 720 363 721
rect 363 720 364 721
rect 365 720 366 721
rect 360 721 366 725
rect 360 725 361 726
rect 362 725 363 726
rect 363 725 364 726
rect 365 725 366 726
rect 400 660 401 661
rect 402 660 403 661
rect 403 660 404 661
rect 405 660 406 661
rect 400 661 406 665
rect 400 665 401 666
rect 402 665 403 666
rect 403 665 404 666
rect 405 665 406 666
rect 640 820 641 821
rect 642 820 643 821
rect 643 820 644 821
rect 645 820 646 821
rect 640 821 646 825
rect 640 825 641 826
rect 642 825 643 826
rect 643 825 644 826
rect 645 825 646 826
rect 240 700 241 701
rect 242 700 243 701
rect 243 700 244 701
rect 245 700 246 701
rect 240 701 246 705
rect 240 705 241 706
rect 242 705 243 706
rect 243 705 244 706
rect 245 705 246 706
rect 620 800 621 801
rect 622 800 623 801
rect 623 800 624 801
rect 625 800 626 801
rect 620 801 626 805
rect 620 805 621 806
rect 622 805 623 806
rect 623 805 624 806
rect 625 805 626 806
rect 260 480 261 481
rect 262 480 263 481
rect 263 480 264 481
rect 265 480 266 481
rect 260 481 266 485
rect 260 485 261 486
rect 262 485 263 486
rect 263 485 264 486
rect 265 485 266 486
rect 740 460 741 461
rect 742 460 743 461
rect 743 460 744 461
rect 745 460 746 461
rect 740 461 746 465
rect 740 465 741 466
rect 742 465 743 466
rect 743 465 744 466
rect 745 465 746 466
rect 680 700 681 701
rect 682 700 683 701
rect 683 700 684 701
rect 685 700 686 701
rect 680 701 686 705
rect 680 705 681 706
rect 682 705 683 706
rect 683 705 684 706
rect 685 705 686 706
rect 520 720 521 721
rect 522 720 523 721
rect 523 720 524 721
rect 525 720 526 721
rect 520 721 526 725
rect 520 725 521 726
rect 522 725 523 726
rect 523 725 524 726
rect 525 725 526 726
rect 600 340 601 341
rect 602 340 603 341
rect 603 340 604 341
rect 605 340 606 341
rect 600 341 606 345
rect 600 345 601 346
rect 602 345 603 346
rect 603 345 604 346
rect 605 345 606 346
rect 440 860 441 861
rect 442 860 443 861
rect 443 860 444 861
rect 445 860 446 861
rect 440 861 446 865
rect 440 865 441 866
rect 442 865 443 866
rect 443 865 444 866
rect 445 865 446 866
rect 560 480 561 481
rect 562 480 563 481
rect 563 480 564 481
rect 565 480 566 481
rect 560 481 566 485
rect 560 485 561 486
rect 562 485 563 486
rect 563 485 564 486
rect 565 485 566 486
rect 680 260 681 261
rect 682 260 683 261
rect 683 260 684 261
rect 685 260 686 261
rect 680 261 686 265
rect 680 265 681 266
rect 682 265 683 266
rect 683 265 684 266
rect 685 265 686 266
rect 480 400 481 401
rect 482 400 483 401
rect 483 400 484 401
rect 485 400 486 401
rect 480 401 486 405
rect 480 405 481 406
rect 482 405 483 406
rect 483 405 484 406
rect 485 405 486 406
rect 720 460 721 461
rect 722 460 723 461
rect 723 460 724 461
rect 725 460 726 461
rect 720 461 726 465
rect 720 465 721 466
rect 722 465 723 466
rect 723 465 724 466
rect 725 465 726 466
rect 380 240 381 241
rect 382 240 383 241
rect 383 240 384 241
rect 385 240 386 241
rect 380 241 386 245
rect 380 245 381 246
rect 382 245 383 246
rect 383 245 384 246
rect 385 245 386 246
rect 440 680 441 681
rect 442 680 443 681
rect 443 680 444 681
rect 445 680 446 681
rect 440 681 446 685
rect 440 685 441 686
rect 442 685 443 686
rect 443 685 444 686
rect 445 685 446 686
rect 400 740 401 741
rect 402 740 403 741
rect 403 740 404 741
rect 405 740 406 741
rect 400 741 406 745
rect 400 745 401 746
rect 402 745 403 746
rect 403 745 404 746
rect 405 745 406 746
rect 640 420 641 421
rect 642 420 643 421
rect 643 420 644 421
rect 645 420 646 421
rect 640 421 646 425
rect 640 425 641 426
rect 642 425 643 426
rect 643 425 644 426
rect 645 425 646 426
rect 280 520 281 521
rect 282 520 283 521
rect 283 520 284 521
rect 285 520 286 521
rect 280 521 286 525
rect 280 525 281 526
rect 282 525 283 526
rect 283 525 284 526
rect 285 525 286 526
rect 700 560 701 561
rect 702 560 703 561
rect 703 560 704 561
rect 705 560 706 561
rect 700 561 706 565
rect 700 565 701 566
rect 702 565 703 566
rect 703 565 704 566
rect 705 565 706 566
rect 340 620 341 621
rect 342 620 343 621
rect 343 620 344 621
rect 345 620 346 621
rect 340 621 346 625
rect 340 625 341 626
rect 342 625 343 626
rect 343 625 344 626
rect 345 625 346 626
rect 520 440 521 441
rect 522 440 523 441
rect 523 440 524 441
rect 525 440 526 441
rect 520 441 526 445
rect 520 445 521 446
rect 522 445 523 446
rect 523 445 524 446
rect 525 445 526 446
rect 540 160 541 161
rect 542 160 543 161
rect 543 160 544 161
rect 545 160 546 161
rect 540 161 546 165
rect 540 165 541 166
rect 542 165 543 166
rect 543 165 544 166
rect 545 165 546 166
rect 440 340 441 341
rect 442 340 443 341
rect 443 340 444 341
rect 445 340 446 341
rect 440 341 446 345
rect 440 345 441 346
rect 442 345 443 346
rect 443 345 444 346
rect 445 345 446 346
rect 800 560 801 561
rect 802 560 803 561
rect 803 560 804 561
rect 805 560 806 561
rect 800 561 806 565
rect 800 565 801 566
rect 802 565 803 566
rect 803 565 804 566
rect 805 565 806 566
rect 480 820 481 821
rect 482 820 483 821
rect 483 820 484 821
rect 485 820 486 821
rect 480 821 486 825
rect 480 825 481 826
rect 482 825 483 826
rect 483 825 484 826
rect 485 825 486 826
rect 240 620 241 621
rect 242 620 243 621
rect 243 620 244 621
rect 245 620 246 621
rect 240 621 246 625
rect 240 625 241 626
rect 242 625 243 626
rect 243 625 244 626
rect 245 625 246 626
rect 320 780 321 781
rect 322 780 323 781
rect 323 780 324 781
rect 325 780 326 781
rect 320 781 326 785
rect 320 785 321 786
rect 322 785 323 786
rect 323 785 324 786
rect 325 785 326 786
rect 360 620 361 621
rect 362 620 363 621
rect 363 620 364 621
rect 365 620 366 621
rect 360 621 366 625
rect 360 625 361 626
rect 362 625 363 626
rect 363 625 364 626
rect 365 625 366 626
rect 700 760 701 761
rect 702 760 703 761
rect 703 760 704 761
rect 705 760 706 761
rect 700 761 706 765
rect 700 765 701 766
rect 702 765 703 766
rect 703 765 704 766
rect 705 765 706 766
rect 420 580 421 581
rect 422 580 423 581
rect 423 580 424 581
rect 425 580 426 581
rect 420 581 426 585
rect 420 585 421 586
rect 422 585 423 586
rect 423 585 424 586
rect 425 585 426 586
rect 680 660 681 661
rect 682 660 683 661
rect 683 660 684 661
rect 685 660 686 661
rect 680 661 686 665
rect 680 665 681 666
rect 682 665 683 666
rect 683 665 684 666
rect 685 665 686 666
rect 320 260 321 261
rect 322 260 323 261
rect 323 260 324 261
rect 325 260 326 261
rect 320 261 326 265
rect 320 265 321 266
rect 322 265 323 266
rect 323 265 324 266
rect 325 265 326 266
rect 800 420 801 421
rect 802 420 803 421
rect 803 420 804 421
rect 805 420 806 421
rect 800 421 806 425
rect 800 425 801 426
rect 802 425 803 426
rect 803 425 804 426
rect 805 425 806 426
rect 320 460 321 461
rect 322 460 323 461
rect 323 460 324 461
rect 325 460 326 461
rect 320 461 326 465
rect 320 465 321 466
rect 322 465 323 466
rect 323 465 324 466
rect 325 465 326 466
rect 700 360 701 361
rect 702 360 703 361
rect 703 360 704 361
rect 705 360 706 361
rect 700 361 706 365
rect 700 365 701 366
rect 702 365 703 366
rect 703 365 704 366
rect 705 365 706 366
rect 600 560 601 561
rect 602 560 603 561
rect 603 560 604 561
rect 605 560 606 561
rect 600 561 606 565
rect 600 565 601 566
rect 602 565 603 566
rect 603 565 604 566
rect 605 565 606 566
rect 240 580 241 581
rect 242 580 243 581
rect 243 580 244 581
rect 245 580 246 581
rect 240 581 246 585
rect 240 585 241 586
rect 242 585 243 586
rect 243 585 244 586
rect 245 585 246 586
rect 740 640 741 641
rect 742 640 743 641
rect 743 640 744 641
rect 745 640 746 641
rect 740 641 746 645
rect 740 645 741 646
rect 742 645 743 646
rect 743 645 744 646
rect 745 645 746 646
rect 740 400 741 401
rect 742 400 743 401
rect 743 400 744 401
rect 745 400 746 401
rect 740 401 746 405
rect 740 405 741 406
rect 742 405 743 406
rect 743 405 744 406
rect 745 405 746 406
rect 660 220 661 221
rect 662 220 663 221
rect 663 220 664 221
rect 665 220 666 221
rect 660 221 666 225
rect 660 225 661 226
rect 662 225 663 226
rect 663 225 664 226
rect 665 225 666 226
rect 100 520 101 521
rect 102 520 103 521
rect 103 520 104 521
rect 105 520 106 521
rect 100 521 106 525
rect 100 525 101 526
rect 102 525 103 526
rect 103 525 104 526
rect 105 525 106 526
rect 360 520 361 521
rect 362 520 363 521
rect 363 520 364 521
rect 365 520 366 521
rect 360 521 366 525
rect 360 525 361 526
rect 362 525 363 526
rect 363 525 364 526
rect 365 525 366 526
rect 420 320 421 321
rect 422 320 423 321
rect 423 320 424 321
rect 425 320 426 321
rect 420 321 426 325
rect 420 325 421 326
rect 422 325 423 326
rect 423 325 424 326
rect 425 325 426 326
rect 500 720 501 721
rect 502 720 503 721
rect 503 720 504 721
rect 505 720 506 721
rect 500 721 506 725
rect 500 725 501 726
rect 502 725 503 726
rect 503 725 504 726
rect 505 725 506 726
rect 740 380 741 381
rect 742 380 743 381
rect 743 380 744 381
rect 745 380 746 381
rect 740 381 746 385
rect 740 385 741 386
rect 742 385 743 386
rect 743 385 744 386
rect 745 385 746 386
rect 220 680 221 681
rect 222 680 223 681
rect 223 680 224 681
rect 225 680 226 681
rect 220 681 226 685
rect 220 685 221 686
rect 222 685 223 686
rect 223 685 224 686
rect 225 685 226 686
rect 420 360 421 361
rect 422 360 423 361
rect 423 360 424 361
rect 425 360 426 361
rect 420 361 426 365
rect 420 365 421 366
rect 422 365 423 366
rect 423 365 424 366
rect 425 365 426 366
rect 260 520 261 521
rect 262 520 263 521
rect 263 520 264 521
rect 265 520 266 521
rect 260 521 266 525
rect 260 525 261 526
rect 262 525 263 526
rect 263 525 264 526
rect 265 525 266 526
rect 780 420 781 421
rect 782 420 783 421
rect 783 420 784 421
rect 785 420 786 421
rect 780 421 786 425
rect 780 425 781 426
rect 782 425 783 426
rect 783 425 784 426
rect 785 425 786 426
rect 380 640 381 641
rect 382 640 383 641
rect 383 640 384 641
rect 385 640 386 641
rect 380 641 386 645
rect 380 645 381 646
rect 382 645 383 646
rect 383 645 384 646
rect 385 645 386 646
rect 520 540 521 541
rect 522 540 523 541
rect 523 540 524 541
rect 525 540 526 541
rect 520 541 526 545
rect 520 545 521 546
rect 522 545 523 546
rect 523 545 524 546
rect 525 545 526 546
rect 720 580 721 581
rect 722 580 723 581
rect 723 580 724 581
rect 725 580 726 581
rect 720 581 726 585
rect 720 585 721 586
rect 722 585 723 586
rect 723 585 724 586
rect 725 585 726 586
rect 440 460 441 461
rect 442 460 443 461
rect 443 460 444 461
rect 445 460 446 461
rect 440 461 446 465
rect 440 465 441 466
rect 442 465 443 466
rect 443 465 444 466
rect 445 465 446 466
rect 660 380 661 381
rect 662 380 663 381
rect 663 380 664 381
rect 665 380 666 381
rect 660 381 666 385
rect 660 385 661 386
rect 662 385 663 386
rect 663 385 664 386
rect 665 385 666 386
rect 420 260 421 261
rect 422 260 423 261
rect 423 260 424 261
rect 425 260 426 261
rect 420 261 426 265
rect 420 265 421 266
rect 422 265 423 266
rect 423 265 424 266
rect 425 265 426 266
rect 520 700 521 701
rect 522 700 523 701
rect 523 700 524 701
rect 525 700 526 701
rect 520 701 526 705
rect 520 705 521 706
rect 522 705 523 706
rect 523 705 524 706
rect 525 705 526 706
rect 680 480 681 481
rect 682 480 683 481
rect 683 480 684 481
rect 685 480 686 481
rect 680 481 686 485
rect 680 485 681 486
rect 682 485 683 486
rect 683 485 684 486
rect 685 485 686 486
rect 680 440 681 441
rect 682 440 683 441
rect 683 440 684 441
rect 685 440 686 441
rect 680 441 686 445
rect 680 445 681 446
rect 682 445 683 446
rect 683 445 684 446
rect 685 445 686 446
rect 360 560 361 561
rect 362 560 363 561
rect 363 560 364 561
rect 365 560 366 561
rect 360 561 366 565
rect 360 565 361 566
rect 362 565 363 566
rect 363 565 364 566
rect 365 565 366 566
rect 600 220 601 221
rect 602 220 603 221
rect 603 220 604 221
rect 605 220 606 221
rect 600 221 606 225
rect 600 225 601 226
rect 602 225 603 226
rect 603 225 604 226
rect 605 225 606 226
rect 520 780 521 781
rect 522 780 523 781
rect 523 780 524 781
rect 525 780 526 781
rect 520 781 526 785
rect 520 785 521 786
rect 522 785 523 786
rect 523 785 524 786
rect 525 785 526 786
rect 260 680 261 681
rect 262 680 263 681
rect 263 680 264 681
rect 265 680 266 681
rect 260 681 266 685
rect 260 685 261 686
rect 262 685 263 686
rect 263 685 264 686
rect 265 685 266 686
rect 540 440 541 441
rect 542 440 543 441
rect 543 440 544 441
rect 545 440 546 441
rect 540 441 546 445
rect 540 445 541 446
rect 542 445 543 446
rect 543 445 544 446
rect 545 445 546 446
rect 320 700 321 701
rect 322 700 323 701
rect 323 700 324 701
rect 325 700 326 701
rect 320 701 326 705
rect 320 705 321 706
rect 322 705 323 706
rect 323 705 324 706
rect 325 705 326 706
rect 760 380 761 381
rect 762 380 763 381
rect 763 380 764 381
rect 765 380 766 381
rect 760 381 766 385
rect 760 385 761 386
rect 762 385 763 386
rect 763 385 764 386
rect 765 385 766 386
rect 420 660 421 661
rect 422 660 423 661
rect 423 660 424 661
rect 425 660 426 661
rect 420 661 426 665
rect 420 665 421 666
rect 422 665 423 666
rect 423 665 424 666
rect 425 665 426 666
rect 220 440 221 441
rect 222 440 223 441
rect 223 440 224 441
rect 225 440 226 441
rect 220 441 226 445
rect 220 445 221 446
rect 222 445 223 446
rect 223 445 224 446
rect 225 445 226 446
rect 360 420 361 421
rect 362 420 363 421
rect 363 420 364 421
rect 365 420 366 421
rect 360 421 366 425
rect 360 425 361 426
rect 362 425 363 426
rect 363 425 364 426
rect 365 425 366 426
rect 780 660 781 661
rect 782 660 783 661
rect 783 660 784 661
rect 785 660 786 661
rect 780 661 786 665
rect 780 665 781 666
rect 782 665 783 666
rect 783 665 784 666
rect 785 665 786 666
rect 460 800 461 801
rect 462 800 463 801
rect 463 800 464 801
rect 465 800 466 801
rect 460 801 466 805
rect 460 805 461 806
rect 462 805 463 806
rect 463 805 464 806
rect 465 805 466 806
rect 720 660 721 661
rect 722 660 723 661
rect 723 660 724 661
rect 725 660 726 661
rect 720 661 726 665
rect 720 665 721 666
rect 722 665 723 666
rect 723 665 724 666
rect 725 665 726 666
rect 560 360 561 361
rect 562 360 563 361
rect 563 360 564 361
rect 565 360 566 361
rect 560 361 566 365
rect 560 365 561 366
rect 562 365 563 366
rect 563 365 564 366
rect 565 365 566 366
rect 600 280 601 281
rect 602 280 603 281
rect 603 280 604 281
rect 605 280 606 281
rect 600 281 606 285
rect 600 285 601 286
rect 602 285 603 286
rect 603 285 604 286
rect 605 285 606 286
rect 380 460 381 461
rect 382 460 383 461
rect 383 460 384 461
rect 385 460 386 461
rect 380 461 386 465
rect 380 465 381 466
rect 382 465 383 466
rect 383 465 384 466
rect 385 465 386 466
rect 580 400 581 401
rect 582 400 583 401
rect 583 400 584 401
rect 585 400 586 401
rect 580 401 586 405
rect 580 405 581 406
rect 582 405 583 406
rect 583 405 584 406
rect 585 405 586 406
rect 520 260 521 261
rect 522 260 523 261
rect 523 260 524 261
rect 525 260 526 261
rect 520 261 526 265
rect 520 265 521 266
rect 522 265 523 266
rect 523 265 524 266
rect 525 265 526 266
rect 620 300 621 301
rect 622 300 623 301
rect 623 300 624 301
rect 625 300 626 301
rect 620 301 626 305
rect 620 305 621 306
rect 622 305 623 306
rect 623 305 624 306
rect 625 305 626 306
rect 280 460 281 461
rect 282 460 283 461
rect 283 460 284 461
rect 285 460 286 461
rect 280 461 286 465
rect 280 465 281 466
rect 282 465 283 466
rect 283 465 284 466
rect 285 465 286 466
rect 300 440 301 441
rect 302 440 303 441
rect 303 440 304 441
rect 305 440 306 441
rect 300 441 306 445
rect 300 445 301 446
rect 302 445 303 446
rect 303 445 304 446
rect 305 445 306 446
rect 500 200 501 201
rect 502 200 503 201
rect 503 200 504 201
rect 505 200 506 201
rect 500 201 506 205
rect 500 205 501 206
rect 502 205 503 206
rect 503 205 504 206
rect 505 205 506 206
rect 140 640 141 641
rect 142 640 143 641
rect 143 640 144 641
rect 145 640 146 641
rect 140 641 146 645
rect 140 645 141 646
rect 142 645 143 646
rect 143 645 144 646
rect 145 645 146 646
rect 640 620 641 621
rect 642 620 643 621
rect 643 620 644 621
rect 645 620 646 621
rect 640 621 646 625
rect 640 625 641 626
rect 642 625 643 626
rect 643 625 644 626
rect 645 625 646 626
rect 400 340 401 341
rect 402 340 403 341
rect 403 340 404 341
rect 405 340 406 341
rect 400 341 406 345
rect 400 345 401 346
rect 402 345 403 346
rect 403 345 404 346
rect 405 345 406 346
rect 880 540 881 541
rect 882 540 883 541
rect 883 540 884 541
rect 885 540 886 541
rect 880 541 886 545
rect 880 545 881 546
rect 882 545 883 546
rect 883 545 884 546
rect 885 545 886 546
rect 760 520 761 521
rect 762 520 763 521
rect 763 520 764 521
rect 765 520 766 521
rect 760 521 766 525
rect 760 525 761 526
rect 762 525 763 526
rect 763 525 764 526
rect 765 525 766 526
rect 420 460 421 461
rect 422 460 423 461
rect 423 460 424 461
rect 425 460 426 461
rect 420 461 426 465
rect 420 465 421 466
rect 422 465 423 466
rect 423 465 424 466
rect 425 465 426 466
rect 480 420 481 421
rect 482 420 483 421
rect 483 420 484 421
rect 485 420 486 421
rect 480 421 486 425
rect 480 425 481 426
rect 482 425 483 426
rect 483 425 484 426
rect 485 425 486 426
rect 520 840 521 841
rect 522 840 523 841
rect 523 840 524 841
rect 525 840 526 841
rect 520 841 526 845
rect 520 845 521 846
rect 522 845 523 846
rect 523 845 524 846
rect 525 845 526 846
rect 540 660 541 661
rect 542 660 543 661
rect 543 660 544 661
rect 545 660 546 661
rect 540 661 546 665
rect 540 665 541 666
rect 542 665 543 666
rect 543 665 544 666
rect 545 665 546 666
rect 460 600 461 601
rect 462 600 463 601
rect 463 600 464 601
rect 465 600 466 601
rect 460 601 466 605
rect 460 605 461 606
rect 462 605 463 606
rect 463 605 464 606
rect 465 605 466 606
rect 460 500 461 501
rect 462 500 463 501
rect 463 500 464 501
rect 465 500 466 501
rect 460 501 466 505
rect 460 505 461 506
rect 462 505 463 506
rect 463 505 464 506
rect 465 505 466 506
rect 780 500 781 501
rect 782 500 783 501
rect 783 500 784 501
rect 785 500 786 501
rect 780 501 786 505
rect 780 505 781 506
rect 782 505 783 506
rect 783 505 784 506
rect 785 505 786 506
rect 340 760 341 761
rect 342 760 343 761
rect 343 760 344 761
rect 345 760 346 761
rect 340 761 346 765
rect 340 765 341 766
rect 342 765 343 766
rect 343 765 344 766
rect 345 765 346 766
rect 260 400 261 401
rect 262 400 263 401
rect 263 400 264 401
rect 265 400 266 401
rect 260 401 266 405
rect 260 405 261 406
rect 262 405 263 406
rect 263 405 264 406
rect 265 405 266 406
rect 440 280 441 281
rect 442 280 443 281
rect 443 280 444 281
rect 445 280 446 281
rect 440 281 446 285
rect 440 285 441 286
rect 442 285 443 286
rect 443 285 444 286
rect 445 285 446 286
rect 680 180 681 181
rect 682 180 683 181
rect 683 180 684 181
rect 685 180 686 181
rect 680 181 686 185
rect 680 185 681 186
rect 682 185 683 186
rect 683 185 684 186
rect 685 185 686 186
rect 220 500 221 501
rect 222 500 223 501
rect 223 500 224 501
rect 225 500 226 501
rect 220 501 226 505
rect 220 505 221 506
rect 222 505 223 506
rect 223 505 224 506
rect 225 505 226 506
rect 620 840 621 841
rect 622 840 623 841
rect 623 840 624 841
rect 625 840 626 841
rect 620 841 626 845
rect 620 845 621 846
rect 622 845 623 846
rect 623 845 624 846
rect 625 845 626 846
rect 540 240 541 241
rect 542 240 543 241
rect 543 240 544 241
rect 545 240 546 241
rect 540 241 546 245
rect 540 245 541 246
rect 542 245 543 246
rect 543 245 544 246
rect 545 245 546 246
rect 360 380 361 381
rect 362 380 363 381
rect 363 380 364 381
rect 365 380 366 381
rect 360 381 366 385
rect 360 385 361 386
rect 362 385 363 386
rect 363 385 364 386
rect 365 385 366 386
rect 720 480 721 481
rect 722 480 723 481
rect 723 480 724 481
rect 725 480 726 481
rect 720 481 726 485
rect 720 485 721 486
rect 722 485 723 486
rect 723 485 724 486
rect 725 485 726 486
rect 280 620 281 621
rect 282 620 283 621
rect 283 620 284 621
rect 285 620 286 621
rect 280 621 286 625
rect 280 625 281 626
rect 282 625 283 626
rect 283 625 284 626
rect 285 625 286 626
rect 240 340 241 341
rect 242 340 243 341
rect 243 340 244 341
rect 245 340 246 341
rect 240 341 246 345
rect 240 345 241 346
rect 242 345 243 346
rect 243 345 244 346
rect 245 345 246 346
rect 360 740 361 741
rect 362 740 363 741
rect 363 740 364 741
rect 365 740 366 741
rect 360 741 366 745
rect 360 745 361 746
rect 362 745 363 746
rect 363 745 364 746
rect 365 745 366 746
rect 380 320 381 321
rect 382 320 383 321
rect 383 320 384 321
rect 385 320 386 321
rect 380 321 386 325
rect 380 325 381 326
rect 382 325 383 326
rect 383 325 384 326
rect 385 325 386 326
rect 380 380 381 381
rect 382 380 383 381
rect 383 380 384 381
rect 385 380 386 381
rect 380 381 386 385
rect 380 385 381 386
rect 382 385 383 386
rect 383 385 384 386
rect 385 385 386 386
rect 200 580 201 581
rect 202 580 203 581
rect 203 580 204 581
rect 205 580 206 581
rect 200 581 206 585
rect 200 585 201 586
rect 202 585 203 586
rect 203 585 204 586
rect 205 585 206 586
rect 400 240 401 241
rect 402 240 403 241
rect 403 240 404 241
rect 405 240 406 241
rect 400 241 406 245
rect 400 245 401 246
rect 402 245 403 246
rect 403 245 404 246
rect 405 245 406 246
rect 240 560 241 561
rect 242 560 243 561
rect 243 560 244 561
rect 245 560 246 561
rect 240 561 246 565
rect 240 565 241 566
rect 242 565 243 566
rect 243 565 244 566
rect 245 565 246 566
rect 720 520 721 521
rect 722 520 723 521
rect 723 520 724 521
rect 725 520 726 521
rect 720 521 726 525
rect 720 525 721 526
rect 722 525 723 526
rect 723 525 724 526
rect 725 525 726 526
rect 660 640 661 641
rect 662 640 663 641
rect 663 640 664 641
rect 665 640 666 641
rect 660 641 666 645
rect 660 645 661 646
rect 662 645 663 646
rect 663 645 664 646
rect 665 645 666 646
rect 300 600 301 601
rect 302 600 303 601
rect 303 600 304 601
rect 305 600 306 601
rect 300 601 306 605
rect 300 605 301 606
rect 302 605 303 606
rect 303 605 304 606
rect 305 605 306 606
rect 500 740 501 741
rect 502 740 503 741
rect 503 740 504 741
rect 505 740 506 741
rect 500 741 506 745
rect 500 745 501 746
rect 502 745 503 746
rect 503 745 504 746
rect 505 745 506 746
rect 600 200 601 201
rect 602 200 603 201
rect 603 200 604 201
rect 605 200 606 201
rect 600 201 606 205
rect 600 205 601 206
rect 602 205 603 206
rect 603 205 604 206
rect 605 205 606 206
rect 580 880 581 881
rect 582 880 583 881
rect 583 880 584 881
rect 585 880 586 881
rect 580 881 586 885
rect 580 885 581 886
rect 582 885 583 886
rect 583 885 584 886
rect 585 885 586 886
rect 180 500 181 501
rect 182 500 183 501
rect 183 500 184 501
rect 185 500 186 501
rect 180 501 186 505
rect 180 505 181 506
rect 182 505 183 506
rect 183 505 184 506
rect 185 505 186 506
rect 580 660 581 661
rect 582 660 583 661
rect 583 660 584 661
rect 585 660 586 661
rect 580 661 586 665
rect 580 665 581 666
rect 582 665 583 666
rect 583 665 584 666
rect 585 665 586 666
rect 660 440 661 441
rect 662 440 663 441
rect 663 440 664 441
rect 665 440 666 441
rect 660 441 666 445
rect 660 445 661 446
rect 662 445 663 446
rect 663 445 664 446
rect 665 445 666 446
rect 520 460 521 461
rect 522 460 523 461
rect 523 460 524 461
rect 525 460 526 461
rect 520 461 526 465
rect 520 465 521 466
rect 522 465 523 466
rect 523 465 524 466
rect 525 465 526 466
rect 460 740 461 741
rect 462 740 463 741
rect 463 740 464 741
rect 465 740 466 741
rect 460 741 466 745
rect 460 745 461 746
rect 462 745 463 746
rect 463 745 464 746
rect 465 745 466 746
rect 440 200 441 201
rect 442 200 443 201
rect 443 200 444 201
rect 445 200 446 201
rect 440 201 446 205
rect 440 205 441 206
rect 442 205 443 206
rect 443 205 444 206
rect 445 205 446 206
rect 860 560 861 561
rect 862 560 863 561
rect 863 560 864 561
rect 865 560 866 561
rect 860 561 866 565
rect 860 565 861 566
rect 862 565 863 566
rect 863 565 864 566
rect 865 565 866 566
rect 300 300 301 301
rect 302 300 303 301
rect 303 300 304 301
rect 305 300 306 301
rect 300 301 306 305
rect 300 305 301 306
rect 302 305 303 306
rect 303 305 304 306
rect 305 305 306 306
rect 300 660 301 661
rect 302 660 303 661
rect 303 660 304 661
rect 305 660 306 661
rect 300 661 306 665
rect 300 665 301 666
rect 302 665 303 666
rect 303 665 304 666
rect 305 665 306 666
rect 760 400 761 401
rect 762 400 763 401
rect 763 400 764 401
rect 765 400 766 401
rect 760 401 766 405
rect 760 405 761 406
rect 762 405 763 406
rect 763 405 764 406
rect 765 405 766 406
rect 340 480 341 481
rect 342 480 343 481
rect 343 480 344 481
rect 345 480 346 481
rect 340 481 346 485
rect 340 485 341 486
rect 342 485 343 486
rect 343 485 344 486
rect 345 485 346 486
rect 480 180 481 181
rect 482 180 483 181
rect 483 180 484 181
rect 485 180 486 181
rect 480 181 486 185
rect 480 185 481 186
rect 482 185 483 186
rect 483 185 484 186
rect 485 185 486 186
rect 240 520 241 521
rect 242 520 243 521
rect 243 520 244 521
rect 245 520 246 521
rect 240 521 246 525
rect 240 525 241 526
rect 242 525 243 526
rect 243 525 244 526
rect 245 525 246 526
rect 640 720 641 721
rect 642 720 643 721
rect 643 720 644 721
rect 645 720 646 721
rect 640 721 646 725
rect 640 725 641 726
rect 642 725 643 726
rect 643 725 644 726
rect 645 725 646 726
rect 440 320 441 321
rect 442 320 443 321
rect 443 320 444 321
rect 445 320 446 321
rect 440 321 446 325
rect 440 325 441 326
rect 442 325 443 326
rect 443 325 444 326
rect 445 325 446 326
rect 800 540 801 541
rect 802 540 803 541
rect 803 540 804 541
rect 805 540 806 541
rect 800 541 806 545
rect 800 545 801 546
rect 802 545 803 546
rect 803 545 804 546
rect 805 545 806 546
rect 340 540 341 541
rect 342 540 343 541
rect 343 540 344 541
rect 345 540 346 541
rect 340 541 346 545
rect 340 545 341 546
rect 342 545 343 546
rect 343 545 344 546
rect 345 545 346 546
rect 540 280 541 281
rect 542 280 543 281
rect 543 280 544 281
rect 545 280 546 281
rect 540 281 546 285
rect 540 285 541 286
rect 542 285 543 286
rect 543 285 544 286
rect 545 285 546 286
rect 700 400 701 401
rect 702 400 703 401
rect 703 400 704 401
rect 705 400 706 401
rect 700 401 706 405
rect 700 405 701 406
rect 702 405 703 406
rect 703 405 704 406
rect 705 405 706 406
rect 540 580 541 581
rect 542 580 543 581
rect 543 580 544 581
rect 545 580 546 581
rect 540 581 546 585
rect 540 585 541 586
rect 542 585 543 586
rect 543 585 544 586
rect 545 585 546 586
rect 320 800 321 801
rect 322 800 323 801
rect 323 800 324 801
rect 325 800 326 801
rect 320 801 326 805
rect 320 805 321 806
rect 322 805 323 806
rect 323 805 324 806
rect 325 805 326 806
rect 340 500 341 501
rect 342 500 343 501
rect 343 500 344 501
rect 345 500 346 501
rect 340 501 346 505
rect 340 505 341 506
rect 342 505 343 506
rect 343 505 344 506
rect 345 505 346 506
rect 540 680 541 681
rect 542 680 543 681
rect 543 680 544 681
rect 545 680 546 681
rect 540 681 546 685
rect 540 685 541 686
rect 542 685 543 686
rect 543 685 544 686
rect 545 685 546 686
rect 560 700 561 701
rect 562 700 563 701
rect 563 700 564 701
rect 565 700 566 701
rect 560 701 566 705
rect 560 705 561 706
rect 562 705 563 706
rect 563 705 564 706
rect 565 705 566 706
rect 720 300 721 301
rect 722 300 723 301
rect 723 300 724 301
rect 725 300 726 301
rect 720 301 726 305
rect 720 305 721 306
rect 722 305 723 306
rect 723 305 724 306
rect 725 305 726 306
rect 560 220 561 221
rect 562 220 563 221
rect 563 220 564 221
rect 565 220 566 221
rect 560 221 566 225
rect 560 225 561 226
rect 562 225 563 226
rect 563 225 564 226
rect 565 225 566 226
rect 420 220 421 221
rect 422 220 423 221
rect 423 220 424 221
rect 425 220 426 221
rect 420 221 426 225
rect 420 225 421 226
rect 422 225 423 226
rect 423 225 424 226
rect 425 225 426 226
rect 520 220 521 221
rect 522 220 523 221
rect 523 220 524 221
rect 525 220 526 221
rect 520 221 526 225
rect 520 225 521 226
rect 522 225 523 226
rect 523 225 524 226
rect 525 225 526 226
rect 280 380 281 381
rect 282 380 283 381
rect 283 380 284 381
rect 285 380 286 381
rect 280 381 286 385
rect 280 385 281 386
rect 282 385 283 386
rect 283 385 284 386
rect 285 385 286 386
rect 760 420 761 421
rect 762 420 763 421
rect 763 420 764 421
rect 765 420 766 421
rect 760 421 766 425
rect 760 425 761 426
rect 762 425 763 426
rect 763 425 764 426
rect 765 425 766 426
rect 500 540 501 541
rect 502 540 503 541
rect 503 540 504 541
rect 505 540 506 541
rect 500 541 506 545
rect 500 545 501 546
rect 502 545 503 546
rect 503 545 504 546
rect 505 545 506 546
rect 440 560 441 561
rect 442 560 443 561
rect 443 560 444 561
rect 445 560 446 561
rect 440 561 446 565
rect 440 565 441 566
rect 442 565 443 566
rect 443 565 444 566
rect 445 565 446 566
rect 520 620 521 621
rect 522 620 523 621
rect 523 620 524 621
rect 525 620 526 621
rect 520 621 526 625
rect 520 625 521 626
rect 522 625 523 626
rect 523 625 524 626
rect 525 625 526 626
rect 120 520 121 521
rect 122 520 123 521
rect 123 520 124 521
rect 125 520 126 521
rect 120 521 126 525
rect 120 525 121 526
rect 122 525 123 526
rect 123 525 124 526
rect 125 525 126 526
rect 600 700 601 701
rect 602 700 603 701
rect 603 700 604 701
rect 605 700 606 701
rect 600 701 606 705
rect 600 705 601 706
rect 602 705 603 706
rect 603 705 604 706
rect 605 705 606 706
rect 880 480 881 481
rect 882 480 883 481
rect 883 480 884 481
rect 885 480 886 481
rect 880 481 886 485
rect 880 485 881 486
rect 882 485 883 486
rect 883 485 884 486
rect 885 485 886 486
rect 640 460 641 461
rect 642 460 643 461
rect 643 460 644 461
rect 645 460 646 461
rect 640 461 646 465
rect 640 465 641 466
rect 642 465 643 466
rect 643 465 644 466
rect 645 465 646 466
rect 500 820 501 821
rect 502 820 503 821
rect 503 820 504 821
rect 505 820 506 821
rect 500 821 506 825
rect 500 825 501 826
rect 502 825 503 826
rect 503 825 504 826
rect 505 825 506 826
rect 500 460 501 461
rect 502 460 503 461
rect 503 460 504 461
rect 505 460 506 461
rect 500 461 506 465
rect 500 465 501 466
rect 502 465 503 466
rect 503 465 504 466
rect 505 465 506 466
rect 300 580 301 581
rect 302 580 303 581
rect 303 580 304 581
rect 305 580 306 581
rect 300 581 306 585
rect 300 585 301 586
rect 302 585 303 586
rect 303 585 304 586
rect 305 585 306 586
rect 640 280 641 281
rect 642 280 643 281
rect 643 280 644 281
rect 645 280 646 281
rect 640 281 646 285
rect 640 285 641 286
rect 642 285 643 286
rect 643 285 644 286
rect 645 285 646 286
rect 400 320 401 321
rect 402 320 403 321
rect 403 320 404 321
rect 405 320 406 321
rect 400 321 406 325
rect 400 325 401 326
rect 402 325 403 326
rect 403 325 404 326
rect 405 325 406 326
rect 280 320 281 321
rect 282 320 283 321
rect 283 320 284 321
rect 285 320 286 321
rect 280 321 286 325
rect 280 325 281 326
rect 282 325 283 326
rect 283 325 284 326
rect 285 325 286 326
rect 800 360 801 361
rect 802 360 803 361
rect 803 360 804 361
rect 805 360 806 361
rect 800 361 806 365
rect 800 365 801 366
rect 802 365 803 366
rect 803 365 804 366
rect 805 365 806 366
rect 620 680 621 681
rect 622 680 623 681
rect 623 680 624 681
rect 625 680 626 681
rect 620 681 626 685
rect 620 685 621 686
rect 622 685 623 686
rect 623 685 624 686
rect 625 685 626 686
rect 520 200 521 201
rect 522 200 523 201
rect 523 200 524 201
rect 525 200 526 201
rect 520 201 526 205
rect 520 205 521 206
rect 522 205 523 206
rect 523 205 524 206
rect 525 205 526 206
rect 840 560 841 561
rect 842 560 843 561
rect 843 560 844 561
rect 845 560 846 561
rect 840 561 846 565
rect 840 565 841 566
rect 842 565 843 566
rect 843 565 844 566
rect 845 565 846 566
rect 440 580 441 581
rect 442 580 443 581
rect 443 580 444 581
rect 445 580 446 581
rect 440 581 446 585
rect 440 585 441 586
rect 442 585 443 586
rect 443 585 444 586
rect 445 585 446 586
rect 500 620 501 621
rect 502 620 503 621
rect 503 620 504 621
rect 505 620 506 621
rect 500 621 506 625
rect 500 625 501 626
rect 502 625 503 626
rect 503 625 504 626
rect 505 625 506 626
rect 500 560 501 561
rect 502 560 503 561
rect 503 560 504 561
rect 505 560 506 561
rect 500 561 506 565
rect 500 565 501 566
rect 502 565 503 566
rect 503 565 504 566
rect 505 565 506 566
rect 280 560 281 561
rect 282 560 283 561
rect 283 560 284 561
rect 285 560 286 561
rect 280 561 286 565
rect 280 565 281 566
rect 282 565 283 566
rect 283 565 284 566
rect 285 565 286 566
rect 480 740 481 741
rect 482 740 483 741
rect 483 740 484 741
rect 485 740 486 741
rect 480 741 486 745
rect 480 745 481 746
rect 482 745 483 746
rect 483 745 484 746
rect 485 745 486 746
rect 640 400 641 401
rect 642 400 643 401
rect 643 400 644 401
rect 645 400 646 401
rect 640 401 646 405
rect 640 405 641 406
rect 642 405 643 406
rect 643 405 644 406
rect 645 405 646 406
rect 580 260 581 261
rect 582 260 583 261
rect 583 260 584 261
rect 585 260 586 261
rect 580 261 586 265
rect 580 265 581 266
rect 582 265 583 266
rect 583 265 584 266
rect 585 265 586 266
rect 220 520 221 521
rect 222 520 223 521
rect 223 520 224 521
rect 225 520 226 521
rect 220 521 226 525
rect 220 525 221 526
rect 222 525 223 526
rect 223 525 224 526
rect 225 525 226 526
rect 400 780 401 781
rect 402 780 403 781
rect 403 780 404 781
rect 405 780 406 781
rect 400 781 406 785
rect 400 785 401 786
rect 402 785 403 786
rect 403 785 404 786
rect 405 785 406 786
rect 500 240 501 241
rect 502 240 503 241
rect 503 240 504 241
rect 505 240 506 241
rect 500 241 506 245
rect 500 245 501 246
rect 502 245 503 246
rect 503 245 504 246
rect 505 245 506 246
rect 720 560 721 561
rect 722 560 723 561
rect 723 560 724 561
rect 725 560 726 561
rect 720 561 726 565
rect 720 565 721 566
rect 722 565 723 566
rect 723 565 724 566
rect 725 565 726 566
rect 420 180 421 181
rect 422 180 423 181
rect 423 180 424 181
rect 425 180 426 181
rect 420 181 426 185
rect 420 185 421 186
rect 422 185 423 186
rect 423 185 424 186
rect 425 185 426 186
rect 240 500 241 501
rect 242 500 243 501
rect 243 500 244 501
rect 245 500 246 501
rect 240 501 246 505
rect 240 505 241 506
rect 242 505 243 506
rect 243 505 244 506
rect 245 505 246 506
rect 580 440 581 441
rect 582 440 583 441
rect 583 440 584 441
rect 585 440 586 441
rect 580 441 586 445
rect 580 445 581 446
rect 582 445 583 446
rect 583 445 584 446
rect 585 445 586 446
rect 780 520 781 521
rect 782 520 783 521
rect 783 520 784 521
rect 785 520 786 521
rect 780 521 786 525
rect 780 525 781 526
rect 782 525 783 526
rect 783 525 784 526
rect 785 525 786 526
rect 680 680 681 681
rect 682 680 683 681
rect 683 680 684 681
rect 685 680 686 681
rect 680 681 686 685
rect 680 685 681 686
rect 682 685 683 686
rect 683 685 684 686
rect 685 685 686 686
rect 260 640 261 641
rect 262 640 263 641
rect 263 640 264 641
rect 265 640 266 641
rect 260 641 266 645
rect 260 645 261 646
rect 262 645 263 646
rect 263 645 264 646
rect 265 645 266 646
rect 860 520 861 521
rect 862 520 863 521
rect 863 520 864 521
rect 865 520 866 521
rect 860 521 866 525
rect 860 525 861 526
rect 862 525 863 526
rect 863 525 864 526
rect 865 525 866 526
rect 540 420 541 421
rect 542 420 543 421
rect 543 420 544 421
rect 545 420 546 421
rect 540 421 546 425
rect 540 425 541 426
rect 542 425 543 426
rect 543 425 544 426
rect 545 425 546 426
rect 520 160 521 161
rect 522 160 523 161
rect 523 160 524 161
rect 525 160 526 161
rect 520 161 526 165
rect 520 165 521 166
rect 522 165 523 166
rect 523 165 524 166
rect 525 165 526 166
rect 560 880 561 881
rect 562 880 563 881
rect 563 880 564 881
rect 565 880 566 881
rect 560 881 566 885
rect 560 885 561 886
rect 562 885 563 886
rect 563 885 564 886
rect 565 885 566 886
rect 320 420 321 421
rect 322 420 323 421
rect 323 420 324 421
rect 325 420 326 421
rect 320 421 326 425
rect 320 425 321 426
rect 322 425 323 426
rect 323 425 324 426
rect 325 425 326 426
rect 540 520 541 521
rect 542 520 543 521
rect 543 520 544 521
rect 545 520 546 521
rect 540 521 546 525
rect 540 525 541 526
rect 542 525 543 526
rect 543 525 544 526
rect 545 525 546 526
rect 580 720 581 721
rect 582 720 583 721
rect 583 720 584 721
rect 585 720 586 721
rect 580 721 586 725
rect 580 725 581 726
rect 582 725 583 726
rect 583 725 584 726
rect 585 725 586 726
rect 200 680 201 681
rect 202 680 203 681
rect 203 680 204 681
rect 205 680 206 681
rect 200 681 206 685
rect 200 685 201 686
rect 202 685 203 686
rect 203 685 204 686
rect 205 685 206 686
rect 360 580 361 581
rect 362 580 363 581
rect 363 580 364 581
rect 365 580 366 581
rect 360 581 366 585
rect 360 585 361 586
rect 362 585 363 586
rect 363 585 364 586
rect 365 585 366 586
rect 620 400 621 401
rect 622 400 623 401
rect 623 400 624 401
rect 625 400 626 401
rect 620 401 626 405
rect 620 405 621 406
rect 622 405 623 406
rect 623 405 624 406
rect 625 405 626 406
rect 560 400 561 401
rect 562 400 563 401
rect 563 400 564 401
rect 565 400 566 401
rect 560 401 566 405
rect 560 405 561 406
rect 562 405 563 406
rect 563 405 564 406
rect 565 405 566 406
rect 560 260 561 261
rect 562 260 563 261
rect 563 260 564 261
rect 565 260 566 261
rect 560 261 566 265
rect 560 265 561 266
rect 562 265 563 266
rect 563 265 564 266
rect 565 265 566 266
rect 760 600 761 601
rect 762 600 763 601
rect 763 600 764 601
rect 765 600 766 601
rect 760 601 766 605
rect 760 605 761 606
rect 762 605 763 606
rect 763 605 764 606
rect 765 605 766 606
rect 480 260 481 261
rect 482 260 483 261
rect 483 260 484 261
rect 485 260 486 261
rect 480 261 486 265
rect 480 265 481 266
rect 482 265 483 266
rect 483 265 484 266
rect 485 265 486 266
rect 620 760 621 761
rect 622 760 623 761
rect 623 760 624 761
rect 625 760 626 761
rect 620 761 626 765
rect 620 765 621 766
rect 622 765 623 766
rect 623 765 624 766
rect 625 765 626 766
rect 760 460 761 461
rect 762 460 763 461
rect 763 460 764 461
rect 765 460 766 461
rect 760 461 766 465
rect 760 465 761 466
rect 762 465 763 466
rect 763 465 764 466
rect 765 465 766 466
rect 620 560 621 561
rect 622 560 623 561
rect 623 560 624 561
rect 625 560 626 561
rect 620 561 626 565
rect 620 565 621 566
rect 622 565 623 566
rect 623 565 624 566
rect 625 565 626 566
rect 780 700 781 701
rect 782 700 783 701
rect 783 700 784 701
rect 785 700 786 701
rect 780 701 786 705
rect 780 705 781 706
rect 782 705 783 706
rect 783 705 784 706
rect 785 705 786 706
rect 580 580 581 581
rect 582 580 583 581
rect 583 580 584 581
rect 585 580 586 581
rect 580 581 586 585
rect 580 585 581 586
rect 582 585 583 586
rect 583 585 584 586
rect 585 585 586 586
rect 460 580 461 581
rect 462 580 463 581
rect 463 580 464 581
rect 465 580 466 581
rect 460 581 466 585
rect 460 585 461 586
rect 462 585 463 586
rect 463 585 464 586
rect 465 585 466 586
rect 580 420 581 421
rect 582 420 583 421
rect 583 420 584 421
rect 585 420 586 421
rect 580 421 586 425
rect 580 425 581 426
rect 582 425 583 426
rect 583 425 584 426
rect 585 425 586 426
rect 660 780 661 781
rect 662 780 663 781
rect 663 780 664 781
rect 665 780 666 781
rect 660 781 666 785
rect 660 785 661 786
rect 662 785 663 786
rect 663 785 664 786
rect 665 785 666 786
rect 820 440 821 441
rect 822 440 823 441
rect 823 440 824 441
rect 825 440 826 441
rect 820 441 826 445
rect 820 445 821 446
rect 822 445 823 446
rect 823 445 824 446
rect 825 445 826 446
rect 500 280 501 281
rect 502 280 503 281
rect 503 280 504 281
rect 505 280 506 281
rect 500 281 506 285
rect 500 285 501 286
rect 502 285 503 286
rect 503 285 504 286
rect 505 285 506 286
rect 560 460 561 461
rect 562 460 563 461
rect 563 460 564 461
rect 565 460 566 461
rect 560 461 566 465
rect 560 465 561 466
rect 562 465 563 466
rect 563 465 564 466
rect 565 465 566 466
rect 160 400 161 401
rect 162 400 163 401
rect 163 400 164 401
rect 165 400 166 401
rect 160 401 166 405
rect 160 405 161 406
rect 162 405 163 406
rect 163 405 164 406
rect 165 405 166 406
rect 580 560 581 561
rect 582 560 583 561
rect 583 560 584 561
rect 585 560 586 561
rect 580 561 586 565
rect 580 565 581 566
rect 582 565 583 566
rect 583 565 584 566
rect 585 565 586 566
rect 580 700 581 701
rect 582 700 583 701
rect 583 700 584 701
rect 585 700 586 701
rect 580 701 586 705
rect 580 705 581 706
rect 582 705 583 706
rect 583 705 584 706
rect 585 705 586 706
rect 820 500 821 501
rect 822 500 823 501
rect 823 500 824 501
rect 825 500 826 501
rect 820 501 826 505
rect 820 505 821 506
rect 822 505 823 506
rect 823 505 824 506
rect 825 505 826 506
rect 720 740 721 741
rect 722 740 723 741
rect 723 740 724 741
rect 725 740 726 741
rect 720 741 726 745
rect 720 745 721 746
rect 722 745 723 746
rect 723 745 724 746
rect 725 745 726 746
rect 440 760 441 761
rect 442 760 443 761
rect 443 760 444 761
rect 445 760 446 761
rect 440 761 446 765
rect 440 765 441 766
rect 442 765 443 766
rect 443 765 444 766
rect 445 765 446 766
rect 760 320 761 321
rect 762 320 763 321
rect 763 320 764 321
rect 765 320 766 321
rect 760 321 766 325
rect 760 325 761 326
rect 762 325 763 326
rect 763 325 764 326
rect 765 325 766 326
rect 340 700 341 701
rect 342 700 343 701
rect 343 700 344 701
rect 345 700 346 701
rect 340 701 346 705
rect 340 705 341 706
rect 342 705 343 706
rect 343 705 344 706
rect 345 705 346 706
rect 720 360 721 361
rect 722 360 723 361
rect 723 360 724 361
rect 725 360 726 361
rect 720 361 726 365
rect 720 365 721 366
rect 722 365 723 366
rect 723 365 724 366
rect 725 365 726 366
rect 700 700 701 701
rect 702 700 703 701
rect 703 700 704 701
rect 705 700 706 701
rect 700 701 706 705
rect 700 705 701 706
rect 702 705 703 706
rect 703 705 704 706
rect 705 705 706 706
rect 520 760 521 761
rect 522 760 523 761
rect 523 760 524 761
rect 525 760 526 761
rect 520 761 526 765
rect 520 765 521 766
rect 522 765 523 766
rect 523 765 524 766
rect 525 765 526 766
rect 520 360 521 361
rect 522 360 523 361
rect 523 360 524 361
rect 525 360 526 361
rect 520 361 526 365
rect 520 365 521 366
rect 522 365 523 366
rect 523 365 524 366
rect 525 365 526 366
rect 420 560 421 561
rect 422 560 423 561
rect 423 560 424 561
rect 425 560 426 561
rect 420 561 426 565
rect 420 565 421 566
rect 422 565 423 566
rect 423 565 424 566
rect 425 565 426 566
rect 160 540 161 541
rect 162 540 163 541
rect 163 540 164 541
rect 165 540 166 541
rect 160 541 166 545
rect 160 545 161 546
rect 162 545 163 546
rect 163 545 164 546
rect 165 545 166 546
rect 340 680 341 681
rect 342 680 343 681
rect 343 680 344 681
rect 345 680 346 681
rect 340 681 346 685
rect 340 685 341 686
rect 342 685 343 686
rect 343 685 344 686
rect 345 685 346 686
rect 680 360 681 361
rect 682 360 683 361
rect 683 360 684 361
rect 685 360 686 361
rect 680 361 686 365
rect 680 365 681 366
rect 682 365 683 366
rect 683 365 684 366
rect 685 365 686 366
rect 220 660 221 661
rect 222 660 223 661
rect 223 660 224 661
rect 225 660 226 661
rect 220 661 226 665
rect 220 665 221 666
rect 222 665 223 666
rect 223 665 224 666
rect 225 665 226 666
rect 140 500 141 501
rect 142 500 143 501
rect 143 500 144 501
rect 145 500 146 501
rect 140 501 146 505
rect 140 505 141 506
rect 142 505 143 506
rect 143 505 144 506
rect 145 505 146 506
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
rect -20 -20 -19 -19
rect -18 -20 -17 -19
rect -17 -20 -16 -19
rect -15 -20 -14 -19
rect -20 -19 -14 -15
rect -20 -15 -19 -14
rect -18 -15 -17 -14
rect -17 -15 -16 -14
rect -15 -15 -14 -14
<< polysilicon >>
rect 361 259 362 261
rect 364 259 365 261
rect 361 265 362 267
rect 364 265 365 267
rect 721 419 722 421
rect 724 419 725 421
rect 721 425 722 427
rect 724 425 725 427
rect 201 379 202 381
rect 204 379 205 381
rect 201 385 202 387
rect 204 385 205 387
rect 741 479 742 481
rect 744 479 745 481
rect 741 485 742 487
rect 744 485 745 487
rect 621 819 622 821
rect 624 819 625 821
rect 621 825 622 827
rect 624 825 625 827
rect 261 539 262 541
rect 264 539 265 541
rect 261 545 262 547
rect 264 545 265 547
rect 381 399 382 401
rect 384 399 385 401
rect 381 405 382 407
rect 384 405 385 407
rect 501 419 502 421
rect 504 419 505 421
rect 501 425 502 427
rect 504 425 505 427
rect 261 359 262 361
rect 264 359 265 361
rect 261 365 262 367
rect 264 365 265 367
rect 261 659 262 661
rect 264 659 265 661
rect 261 665 262 667
rect 264 665 265 667
rect 761 659 762 661
rect 764 659 765 661
rect 761 665 762 667
rect 764 665 765 667
rect 381 659 382 661
rect 384 659 385 661
rect 381 665 382 667
rect 384 665 385 667
rect 481 799 482 801
rect 484 799 485 801
rect 481 805 482 807
rect 484 805 485 807
rect 741 679 742 681
rect 744 679 745 681
rect 741 685 742 687
rect 744 685 745 687
rect 181 479 182 481
rect 184 479 185 481
rect 181 485 182 487
rect 184 485 185 487
rect 601 619 602 621
rect 604 619 605 621
rect 601 625 602 627
rect 604 625 605 627
rect 861 539 862 541
rect 864 539 865 541
rect 861 545 862 547
rect 864 545 865 547
rect 561 579 562 581
rect 564 579 565 581
rect 561 585 562 587
rect 564 585 565 587
rect 661 619 662 621
rect 664 619 665 621
rect 661 625 662 627
rect 664 625 665 627
rect 321 379 322 381
rect 324 379 325 381
rect 321 385 322 387
rect 324 385 325 387
rect 581 799 582 801
rect 584 799 585 801
rect 581 805 582 807
rect 584 805 585 807
rect 201 439 202 441
rect 204 439 205 441
rect 201 445 202 447
rect 204 445 205 447
rect 321 579 322 581
rect 324 579 325 581
rect 321 585 322 587
rect 324 585 325 587
rect 221 359 222 361
rect 224 359 225 361
rect 221 365 222 367
rect 224 365 225 367
rect 261 339 262 341
rect 264 339 265 341
rect 261 345 262 347
rect 264 345 265 347
rect 641 559 642 561
rect 644 559 645 561
rect 641 565 642 567
rect 644 565 645 567
rect 161 439 162 441
rect 164 439 165 441
rect 161 445 162 447
rect 164 445 165 447
rect 621 719 622 721
rect 624 719 625 721
rect 621 725 622 727
rect 624 725 625 727
rect 461 719 462 721
rect 464 719 465 721
rect 461 725 462 727
rect 464 725 465 727
rect 481 659 482 661
rect 484 659 485 661
rect 481 665 482 667
rect 484 665 485 667
rect 601 459 602 461
rect 604 459 605 461
rect 601 465 602 467
rect 604 465 605 467
rect 381 479 382 481
rect 384 479 385 481
rect 381 485 382 487
rect 384 485 385 487
rect 721 679 722 681
rect 724 679 725 681
rect 721 685 722 687
rect 724 685 725 687
rect 541 459 542 461
rect 544 459 545 461
rect 541 465 542 467
rect 544 465 545 467
rect 621 499 622 501
rect 624 499 625 501
rect 621 505 622 507
rect 624 505 625 507
rect 381 279 382 281
rect 384 279 385 281
rect 381 285 382 287
rect 384 285 385 287
rect 821 659 822 661
rect 824 659 825 661
rect 821 665 822 667
rect 824 665 825 667
rect 121 499 122 501
rect 124 499 125 501
rect 121 505 122 507
rect 124 505 125 507
rect 501 799 502 801
rect 504 799 505 801
rect 501 805 502 807
rect 504 805 505 807
rect 641 299 642 301
rect 644 299 645 301
rect 641 305 642 307
rect 644 305 645 307
rect 801 459 802 461
rect 804 459 805 461
rect 801 465 802 467
rect 804 465 805 467
rect 481 279 482 281
rect 484 279 485 281
rect 481 285 482 287
rect 484 285 485 287
rect 741 699 742 701
rect 744 699 745 701
rect 741 705 742 707
rect 744 705 745 707
rect 801 379 802 381
rect 804 379 805 381
rect 801 385 802 387
rect 804 385 805 387
rect 421 679 422 681
rect 424 679 425 681
rect 421 685 422 687
rect 424 685 425 687
rect 441 179 442 181
rect 444 179 445 181
rect 441 185 442 187
rect 444 185 445 187
rect 501 839 502 841
rect 504 839 505 841
rect 501 845 502 847
rect 504 845 505 847
rect 541 639 542 641
rect 544 639 545 641
rect 541 645 542 647
rect 544 645 545 647
rect 621 259 622 261
rect 624 259 625 261
rect 621 265 622 267
rect 624 265 625 267
rect 481 859 482 861
rect 484 859 485 861
rect 481 865 482 867
rect 484 865 485 867
rect 441 799 442 801
rect 444 799 445 801
rect 441 805 442 807
rect 444 805 445 807
rect 821 459 822 461
rect 824 459 825 461
rect 821 465 822 467
rect 824 465 825 467
rect 601 739 602 741
rect 604 739 605 741
rect 601 745 602 747
rect 604 745 605 747
rect 461 679 462 681
rect 464 679 465 681
rect 461 685 462 687
rect 464 685 465 687
rect 221 479 222 481
rect 224 479 225 481
rect 221 485 222 487
rect 224 485 225 487
rect 661 539 662 541
rect 664 539 665 541
rect 661 545 662 547
rect 664 545 665 547
rect 341 719 342 721
rect 344 719 345 721
rect 341 725 342 727
rect 344 725 345 727
rect 441 879 442 881
rect 444 879 445 881
rect 441 885 442 887
rect 444 885 445 887
rect 401 799 402 801
rect 404 799 405 801
rect 401 805 402 807
rect 404 805 405 807
rect 141 579 142 581
rect 144 579 145 581
rect 141 585 142 587
rect 144 585 145 587
rect 181 579 182 581
rect 184 579 185 581
rect 181 585 182 587
rect 184 585 185 587
rect 721 719 722 721
rect 724 719 725 721
rect 721 725 722 727
rect 724 725 725 727
rect 321 479 322 481
rect 324 479 325 481
rect 321 485 322 487
rect 324 485 325 487
rect 621 619 622 621
rect 624 619 625 621
rect 621 625 622 627
rect 624 625 625 627
rect 561 799 562 801
rect 564 799 565 801
rect 561 805 562 807
rect 564 805 565 807
rect 281 759 282 761
rect 284 759 285 761
rect 281 765 282 767
rect 284 765 285 767
rect 801 679 802 681
rect 804 679 805 681
rect 801 685 802 687
rect 804 685 805 687
rect 541 559 542 561
rect 544 559 545 561
rect 541 565 542 567
rect 544 565 545 567
rect 441 499 442 501
rect 444 499 445 501
rect 441 505 442 507
rect 444 505 445 507
rect 781 379 782 381
rect 784 379 785 381
rect 781 385 782 387
rect 784 385 785 387
rect 801 599 802 601
rect 804 599 805 601
rect 801 605 802 607
rect 804 605 805 607
rect 641 699 642 701
rect 644 699 645 701
rect 641 705 642 707
rect 644 705 645 707
rect 501 759 502 761
rect 504 759 505 761
rect 501 765 502 767
rect 504 765 505 767
rect 321 359 322 361
rect 324 359 325 361
rect 321 365 322 367
rect 324 365 325 367
rect 161 559 162 561
rect 164 559 165 561
rect 161 565 162 567
rect 164 565 165 567
rect 421 379 422 381
rect 424 379 425 381
rect 421 385 422 387
rect 424 385 425 387
rect 141 619 142 621
rect 144 619 145 621
rect 141 625 142 627
rect 144 625 145 627
rect 681 579 682 581
rect 684 579 685 581
rect 681 585 682 587
rect 684 585 685 587
rect 781 619 782 621
rect 784 619 785 621
rect 781 625 782 627
rect 784 625 785 627
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect 321 619 322 621
rect 324 619 325 621
rect 321 625 322 627
rect 324 625 325 627
rect 721 439 722 441
rect 724 439 725 441
rect 721 445 722 447
rect 724 445 725 447
rect 481 579 482 581
rect 484 579 485 581
rect 481 585 482 587
rect 484 585 485 587
rect 341 739 342 741
rect 344 739 345 741
rect 341 745 342 747
rect 344 745 345 747
rect 181 639 182 641
rect 184 639 185 641
rect 181 645 182 647
rect 184 645 185 647
rect 801 439 802 441
rect 804 439 805 441
rect 801 445 802 447
rect 804 445 805 447
rect 661 319 662 321
rect 664 319 665 321
rect 661 325 662 327
rect 664 325 665 327
rect 261 739 262 741
rect 264 739 265 741
rect 261 745 262 747
rect 264 745 265 747
rect 381 199 382 201
rect 384 199 385 201
rect 381 205 382 207
rect 384 205 385 207
rect 621 379 622 381
rect 624 379 625 381
rect 621 385 622 387
rect 624 385 625 387
rect 641 799 642 801
rect 644 799 645 801
rect 641 805 642 807
rect 644 805 645 807
rect 481 159 482 161
rect 484 159 485 161
rect 481 165 482 167
rect 484 165 485 167
rect 261 719 262 721
rect 264 719 265 721
rect 261 725 262 727
rect 264 725 265 727
rect 581 479 582 481
rect 584 479 585 481
rect 581 485 582 487
rect 584 485 585 487
rect 441 779 442 781
rect 444 779 445 781
rect 441 785 442 787
rect 444 785 445 787
rect 861 499 862 501
rect 864 499 865 501
rect 861 505 862 507
rect 864 505 865 507
rect 841 399 842 401
rect 844 399 845 401
rect 841 405 842 407
rect 844 405 845 407
rect 321 599 322 601
rect 324 599 325 601
rect 321 605 322 607
rect 324 605 325 607
rect 521 819 522 821
rect 524 819 525 821
rect 521 825 522 827
rect 524 825 525 827
rect 521 859 522 861
rect 524 859 525 861
rect 521 865 522 867
rect 524 865 525 867
rect 481 639 482 641
rect 484 639 485 641
rect 481 645 482 647
rect 484 645 485 647
rect 721 499 722 501
rect 724 499 725 501
rect 721 505 722 507
rect 724 505 725 507
rect 661 199 662 201
rect 664 199 665 201
rect 661 205 662 207
rect 664 205 665 207
rect 401 419 402 421
rect 404 419 405 421
rect 401 425 402 427
rect 404 425 405 427
rect 401 819 402 821
rect 404 819 405 821
rect 401 825 402 827
rect 404 825 405 827
rect 741 299 742 301
rect 744 299 745 301
rect 741 305 742 307
rect 744 305 745 307
rect 461 619 462 621
rect 464 619 465 621
rect 461 625 462 627
rect 464 625 465 627
rect 621 699 622 701
rect 624 699 625 701
rect 621 705 622 707
rect 624 705 625 707
rect 161 579 162 581
rect 164 579 165 581
rect 161 585 162 587
rect 164 585 165 587
rect 461 659 462 661
rect 464 659 465 661
rect 461 665 462 667
rect 464 665 465 667
rect 261 379 262 381
rect 264 379 265 381
rect 261 385 262 387
rect 264 385 265 387
rect 561 639 562 641
rect 564 639 565 641
rect 561 645 562 647
rect 564 645 565 647
rect 341 439 342 441
rect 344 439 345 441
rect 341 445 342 447
rect 344 445 345 447
rect 281 299 282 301
rect 284 299 285 301
rect 281 305 282 307
rect 284 305 285 307
rect 401 259 402 261
rect 404 259 405 261
rect 401 265 402 267
rect 404 265 405 267
rect 501 859 502 861
rect 504 859 505 861
rect 501 865 502 867
rect 504 865 505 867
rect 401 219 402 221
rect 404 219 405 221
rect 401 225 402 227
rect 404 225 405 227
rect 361 219 362 221
rect 364 219 365 221
rect 361 225 362 227
rect 364 225 365 227
rect 761 479 762 481
rect 764 479 765 481
rect 761 485 762 487
rect 764 485 765 487
rect 641 499 642 501
rect 644 499 645 501
rect 641 505 642 507
rect 644 505 645 507
rect 521 579 522 581
rect 524 579 525 581
rect 521 585 522 587
rect 524 585 525 587
rect 381 519 382 521
rect 384 519 385 521
rect 381 525 382 527
rect 384 525 385 527
rect 461 439 462 441
rect 464 439 465 441
rect 461 445 462 447
rect 464 445 465 447
rect 781 359 782 361
rect 784 359 785 361
rect 781 365 782 367
rect 784 365 785 367
rect 541 899 542 901
rect 544 899 545 901
rect 541 905 542 907
rect 544 905 545 907
rect 361 799 362 801
rect 364 799 365 801
rect 361 805 362 807
rect 364 805 365 807
rect 181 539 182 541
rect 184 539 185 541
rect 181 545 182 547
rect 184 545 185 547
rect 261 499 262 501
rect 264 499 265 501
rect 261 505 262 507
rect 264 505 265 507
rect 381 719 382 721
rect 384 719 385 721
rect 381 725 382 727
rect 384 725 385 727
rect 481 299 482 301
rect 484 299 485 301
rect 481 305 482 307
rect 484 305 485 307
rect 301 379 302 381
rect 304 379 305 381
rect 301 385 302 387
rect 304 385 305 387
rect 421 199 422 201
rect 424 199 425 201
rect 421 205 422 207
rect 424 205 425 207
rect 581 199 582 201
rect 584 199 585 201
rect 581 205 582 207
rect 584 205 585 207
rect 561 659 562 661
rect 564 659 565 661
rect 561 665 562 667
rect 564 665 565 667
rect 641 839 642 841
rect 644 839 645 841
rect 641 845 642 847
rect 644 845 645 847
rect 421 599 422 601
rect 424 599 425 601
rect 421 605 422 607
rect 424 605 425 607
rect 281 499 282 501
rect 284 499 285 501
rect 281 505 282 507
rect 284 505 285 507
rect 421 399 422 401
rect 424 399 425 401
rect 421 405 422 407
rect 424 405 425 407
rect 681 399 682 401
rect 684 399 685 401
rect 681 405 682 407
rect 684 405 685 407
rect 241 379 242 381
rect 244 379 245 381
rect 241 385 242 387
rect 244 385 245 387
rect 321 639 322 641
rect 324 639 325 641
rect 321 645 322 647
rect 324 645 325 647
rect 321 339 322 341
rect 324 339 325 341
rect 321 345 322 347
rect 324 345 325 347
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect 401 539 402 541
rect 404 539 405 541
rect 401 545 402 547
rect 404 545 405 547
rect 301 479 302 481
rect 304 479 305 481
rect 301 485 302 487
rect 304 485 305 487
rect 421 339 422 341
rect 424 339 425 341
rect 421 345 422 347
rect 424 345 425 347
rect 821 519 822 521
rect 824 519 825 521
rect 821 525 822 527
rect 824 525 825 527
rect 201 659 202 661
rect 204 659 205 661
rect 201 665 202 667
rect 204 665 205 667
rect 601 419 602 421
rect 604 419 605 421
rect 601 425 602 427
rect 604 425 605 427
rect 821 579 822 581
rect 824 579 825 581
rect 821 585 822 587
rect 824 585 825 587
rect 361 339 362 341
rect 364 339 365 341
rect 361 345 362 347
rect 364 345 365 347
rect 641 539 642 541
rect 644 539 645 541
rect 641 545 642 547
rect 644 545 645 547
rect 641 339 642 341
rect 644 339 645 341
rect 641 345 642 347
rect 644 345 645 347
rect 481 459 482 461
rect 484 459 485 461
rect 481 465 482 467
rect 484 465 485 467
rect 481 339 482 341
rect 484 339 485 341
rect 481 345 482 347
rect 484 345 485 347
rect 361 439 362 441
rect 364 439 365 441
rect 361 445 362 447
rect 364 445 365 447
rect 661 339 662 341
rect 664 339 665 341
rect 661 345 662 347
rect 664 345 665 347
rect 281 739 282 741
rect 284 739 285 741
rect 281 745 282 747
rect 284 745 285 747
rect 701 499 702 501
rect 704 499 705 501
rect 701 505 702 507
rect 704 505 705 507
rect 261 319 262 321
rect 264 319 265 321
rect 261 325 262 327
rect 264 325 265 327
rect 381 339 382 341
rect 384 339 385 341
rect 381 345 382 347
rect 384 345 385 347
rect 701 539 702 541
rect 704 539 705 541
rect 701 545 702 547
rect 704 545 705 547
rect 881 519 882 521
rect 884 519 885 521
rect 881 525 882 527
rect 884 525 885 527
rect 841 539 842 541
rect 844 539 845 541
rect 841 545 842 547
rect 844 545 845 547
rect 621 779 622 781
rect 624 779 625 781
rect 621 785 622 787
rect 624 785 625 787
rect 321 539 322 541
rect 324 539 325 541
rect 321 545 322 547
rect 324 545 325 547
rect 761 699 762 701
rect 764 699 765 701
rect 761 705 762 707
rect 764 705 765 707
rect 361 779 362 781
rect 364 779 365 781
rect 361 785 362 787
rect 364 785 365 787
rect 421 819 422 821
rect 424 819 425 821
rect 421 825 422 827
rect 424 825 425 827
rect 741 719 742 721
rect 744 719 745 721
rect 741 725 742 727
rect 744 725 745 727
rect 681 599 682 601
rect 684 599 685 601
rect 681 605 682 607
rect 684 605 685 607
rect 641 219 642 221
rect 644 219 645 221
rect 641 225 642 227
rect 644 225 645 227
rect 641 319 642 321
rect 644 319 645 321
rect 641 325 642 327
rect 644 325 645 327
rect 781 639 782 641
rect 784 639 785 641
rect 781 645 782 647
rect 784 645 785 647
rect 801 619 802 621
rect 804 619 805 621
rect 801 625 802 627
rect 804 625 805 627
rect 461 219 462 221
rect 464 219 465 221
rect 461 225 462 227
rect 464 225 465 227
rect 501 519 502 521
rect 504 519 505 521
rect 501 525 502 527
rect 504 525 505 527
rect 441 299 442 301
rect 444 299 445 301
rect 441 305 442 307
rect 444 305 445 307
rect 101 459 102 461
rect 104 459 105 461
rect 101 465 102 467
rect 104 465 105 467
rect 181 519 182 521
rect 184 519 185 521
rect 181 525 182 527
rect 184 525 185 527
rect 261 559 262 561
rect 264 559 265 561
rect 261 565 262 567
rect 264 565 265 567
rect 601 399 602 401
rect 604 399 605 401
rect 601 405 602 407
rect 604 405 605 407
rect 521 659 522 661
rect 524 659 525 661
rect 521 665 522 667
rect 524 665 525 667
rect 141 519 142 521
rect 144 519 145 521
rect 141 525 142 527
rect 144 525 145 527
rect 801 399 802 401
rect 804 399 805 401
rect 801 405 802 407
rect 804 405 805 407
rect 581 819 582 821
rect 584 819 585 821
rect 581 825 582 827
rect 584 825 585 827
rect 561 539 562 541
rect 564 539 565 541
rect 561 545 562 547
rect 564 545 565 547
rect 201 499 202 501
rect 204 499 205 501
rect 201 505 202 507
rect 204 505 205 507
rect 701 339 702 341
rect 704 339 705 341
rect 701 345 702 347
rect 704 345 705 347
rect 561 419 562 421
rect 564 419 565 421
rect 561 425 562 427
rect 564 425 565 427
rect 141 599 142 601
rect 144 599 145 601
rect 141 605 142 607
rect 144 605 145 607
rect 501 379 502 381
rect 504 379 505 381
rect 501 385 502 387
rect 504 385 505 387
rect 601 799 602 801
rect 604 799 605 801
rect 601 805 602 807
rect 604 805 605 807
rect 441 619 442 621
rect 444 619 445 621
rect 441 625 442 627
rect 444 625 445 627
rect 201 539 202 541
rect 204 539 205 541
rect 201 545 202 547
rect 204 545 205 547
rect 161 419 162 421
rect 164 419 165 421
rect 161 425 162 427
rect 164 425 165 427
rect 561 159 562 161
rect 564 159 565 161
rect 561 165 562 167
rect 564 165 565 167
rect 381 759 382 761
rect 384 759 385 761
rect 381 765 382 767
rect 384 765 385 767
rect 901 559 902 561
rect 904 559 905 561
rect 901 565 902 567
rect 904 565 905 567
rect 281 599 282 601
rect 284 599 285 601
rect 281 605 282 607
rect 284 605 285 607
rect 521 519 522 521
rect 524 519 525 521
rect 521 525 522 527
rect 524 525 525 527
rect 521 419 522 421
rect 524 419 525 421
rect 521 425 522 427
rect 524 425 525 427
rect 341 259 342 261
rect 344 259 345 261
rect 341 265 342 267
rect 344 265 345 267
rect 201 519 202 521
rect 204 519 205 521
rect 201 525 202 527
rect 204 525 205 527
rect 761 499 762 501
rect 764 499 765 501
rect 761 505 762 507
rect 764 505 765 507
rect 881 499 882 501
rect 884 499 885 501
rect 881 505 882 507
rect 884 505 885 507
rect 361 759 362 761
rect 364 759 365 761
rect 361 765 362 767
rect 364 765 365 767
rect 581 779 582 781
rect 584 779 585 781
rect 581 785 582 787
rect 584 785 585 787
rect 621 179 622 181
rect 624 179 625 181
rect 621 185 622 187
rect 624 185 625 187
rect 341 399 342 401
rect 344 399 345 401
rect 341 405 342 407
rect 344 405 345 407
rect 441 539 442 541
rect 444 539 445 541
rect 441 545 442 547
rect 444 545 445 547
rect 821 599 822 601
rect 824 599 825 601
rect 821 605 822 607
rect 824 605 825 607
rect 361 279 362 281
rect 364 279 365 281
rect 361 285 362 287
rect 364 285 365 287
rect 541 499 542 501
rect 544 499 545 501
rect 541 505 542 507
rect 544 505 545 507
rect 541 179 542 181
rect 544 179 545 181
rect 541 185 542 187
rect 544 185 545 187
rect 401 759 402 761
rect 404 759 405 761
rect 401 765 402 767
rect 404 765 405 767
rect 701 299 702 301
rect 704 299 705 301
rect 701 305 702 307
rect 704 305 705 307
rect 281 539 282 541
rect 284 539 285 541
rect 281 545 282 547
rect 284 545 285 547
rect 781 679 782 681
rect 784 679 785 681
rect 781 685 782 687
rect 784 685 785 687
rect 181 659 182 661
rect 184 659 185 661
rect 181 665 182 667
rect 184 665 185 667
rect 441 239 442 241
rect 444 239 445 241
rect 441 245 442 247
rect 444 245 445 247
rect 341 819 342 821
rect 344 819 345 821
rect 341 825 342 827
rect 344 825 345 827
rect 581 319 582 321
rect 584 319 585 321
rect 581 325 582 327
rect 584 325 585 327
rect 321 719 322 721
rect 324 719 325 721
rect 321 725 322 727
rect 324 725 325 727
rect 501 579 502 581
rect 504 579 505 581
rect 501 585 502 587
rect 504 585 505 587
rect 541 139 542 141
rect 544 139 545 141
rect 541 145 542 147
rect 544 145 545 147
rect 401 559 402 561
rect 404 559 405 561
rect 401 565 402 567
rect 404 565 405 567
rect 661 499 662 501
rect 664 499 665 501
rect 661 505 662 507
rect 664 505 665 507
rect 201 619 202 621
rect 204 619 205 621
rect 201 625 202 627
rect 204 625 205 627
rect 581 759 582 761
rect 584 759 585 761
rect 581 765 582 767
rect 584 765 585 767
rect 121 439 122 441
rect 124 439 125 441
rect 121 445 122 447
rect 124 445 125 447
rect 481 839 482 841
rect 484 839 485 841
rect 481 845 482 847
rect 484 845 485 847
rect 481 759 482 761
rect 484 759 485 761
rect 481 765 482 767
rect 484 765 485 767
rect 301 419 302 421
rect 304 419 305 421
rect 301 425 302 427
rect 304 425 305 427
rect 821 639 822 641
rect 824 639 825 641
rect 821 645 822 647
rect 824 645 825 647
rect 521 559 522 561
rect 524 559 525 561
rect 521 565 522 567
rect 524 565 525 567
rect 501 879 502 881
rect 504 879 505 881
rect 501 885 502 887
rect 504 885 505 887
rect 321 499 322 501
rect 324 499 325 501
rect 321 505 322 507
rect 324 505 325 507
rect 881 459 882 461
rect 884 459 885 461
rect 881 465 882 467
rect 884 465 885 467
rect 581 219 582 221
rect 584 219 585 221
rect 581 225 582 227
rect 584 225 585 227
rect 801 639 802 641
rect 804 639 805 641
rect 801 645 802 647
rect 804 645 805 647
rect 161 519 162 521
rect 164 519 165 521
rect 161 525 162 527
rect 164 525 165 527
rect 641 579 642 581
rect 644 579 645 581
rect 641 585 642 587
rect 644 585 645 587
rect 541 319 542 321
rect 544 319 545 321
rect 541 325 542 327
rect 544 325 545 327
rect 281 439 282 441
rect 284 439 285 441
rect 281 445 282 447
rect 284 445 285 447
rect 601 839 602 841
rect 604 839 605 841
rect 601 845 602 847
rect 604 845 605 847
rect 801 499 802 501
rect 804 499 805 501
rect 801 505 802 507
rect 804 505 805 507
rect 301 719 302 721
rect 304 719 305 721
rect 301 725 302 727
rect 304 725 305 727
rect 681 519 682 521
rect 684 519 685 521
rect 681 525 682 527
rect 684 525 685 527
rect 421 839 422 841
rect 424 839 425 841
rect 421 845 422 847
rect 424 845 425 847
rect 401 439 402 441
rect 404 439 405 441
rect 401 445 402 447
rect 404 445 405 447
rect 441 359 442 361
rect 444 359 445 361
rect 441 365 442 367
rect 444 365 445 367
rect 841 459 842 461
rect 844 459 845 461
rect 841 465 842 467
rect 844 465 845 467
rect 301 739 302 741
rect 304 739 305 741
rect 301 745 302 747
rect 304 745 305 747
rect 281 719 282 721
rect 284 719 285 721
rect 281 725 282 727
rect 284 725 285 727
rect 381 599 382 601
rect 384 599 385 601
rect 381 605 382 607
rect 384 605 385 607
rect 601 819 602 821
rect 604 819 605 821
rect 601 825 602 827
rect 604 825 605 827
rect 481 319 482 321
rect 484 319 485 321
rect 481 325 482 327
rect 484 325 485 327
rect 741 439 742 441
rect 744 439 745 441
rect 741 445 742 447
rect 744 445 745 447
rect 481 539 482 541
rect 484 539 485 541
rect 481 545 482 547
rect 484 545 485 547
rect 541 839 542 841
rect 544 839 545 841
rect 541 845 542 847
rect 544 845 545 847
rect 441 839 442 841
rect 444 839 445 841
rect 441 845 442 847
rect 444 845 445 847
rect 461 859 462 861
rect 464 859 465 861
rect 461 865 462 867
rect 464 865 465 867
rect 301 699 302 701
rect 304 699 305 701
rect 301 705 302 707
rect 304 705 305 707
rect 461 519 462 521
rect 464 519 465 521
rect 461 525 462 527
rect 464 525 465 527
rect 421 799 422 801
rect 424 799 425 801
rect 421 805 422 807
rect 424 805 425 807
rect 521 599 522 601
rect 524 599 525 601
rect 521 605 522 607
rect 524 605 525 607
rect 761 719 762 721
rect 764 719 765 721
rect 761 725 762 727
rect 764 725 765 727
rect 341 559 342 561
rect 344 559 345 561
rect 341 565 342 567
rect 344 565 345 567
rect 501 179 502 181
rect 504 179 505 181
rect 501 185 502 187
rect 504 185 505 187
rect 441 379 442 381
rect 444 379 445 381
rect 441 385 442 387
rect 444 385 445 387
rect 281 339 282 341
rect 284 339 285 341
rect 281 345 282 347
rect 284 345 285 347
rect 221 559 222 561
rect 224 559 225 561
rect 221 565 222 567
rect 224 565 225 567
rect 841 439 842 441
rect 844 439 845 441
rect 841 445 842 447
rect 844 445 845 447
rect 241 679 242 681
rect 244 679 245 681
rect 241 685 242 687
rect 244 685 245 687
rect 501 599 502 601
rect 504 599 505 601
rect 501 605 502 607
rect 504 605 505 607
rect 741 739 742 741
rect 744 739 745 741
rect 741 745 742 747
rect 744 745 745 747
rect 201 359 202 361
rect 204 359 205 361
rect 201 365 202 367
rect 204 365 205 367
rect 161 619 162 621
rect 164 619 165 621
rect 161 625 162 627
rect 164 625 165 627
rect 281 579 282 581
rect 284 579 285 581
rect 281 585 282 587
rect 284 585 285 587
rect 741 599 742 601
rect 744 599 745 601
rect 741 605 742 607
rect 744 605 745 607
rect 461 839 462 841
rect 464 839 465 841
rect 461 845 462 847
rect 464 845 465 847
rect 681 379 682 381
rect 684 379 685 381
rect 681 385 682 387
rect 684 385 685 387
rect 241 439 242 441
rect 244 439 245 441
rect 241 445 242 447
rect 244 445 245 447
rect 641 779 642 781
rect 644 779 645 781
rect 641 785 642 787
rect 644 785 645 787
rect 461 339 462 341
rect 464 339 465 341
rect 461 345 462 347
rect 464 345 465 347
rect 741 659 742 661
rect 744 659 745 661
rect 741 665 742 667
rect 744 665 745 667
rect 361 599 362 601
rect 364 599 365 601
rect 361 605 362 607
rect 364 605 365 607
rect 421 479 422 481
rect 424 479 425 481
rect 421 485 422 487
rect 424 485 425 487
rect 701 659 702 661
rect 704 659 705 661
rect 701 665 702 667
rect 704 665 705 667
rect 341 319 342 321
rect 344 319 345 321
rect 341 325 342 327
rect 344 325 345 327
rect 541 539 542 541
rect 544 539 545 541
rect 541 545 542 547
rect 544 545 545 547
rect 221 459 222 461
rect 224 459 225 461
rect 221 465 222 467
rect 224 465 225 467
rect 861 459 862 461
rect 864 459 865 461
rect 861 465 862 467
rect 864 465 865 467
rect 561 739 562 741
rect 564 739 565 741
rect 561 745 562 747
rect 564 745 565 747
rect 161 599 162 601
rect 164 599 165 601
rect 161 605 162 607
rect 164 605 165 607
rect 641 259 642 261
rect 644 259 645 261
rect 641 265 642 267
rect 644 265 645 267
rect 721 259 722 261
rect 724 259 725 261
rect 721 265 722 267
rect 724 265 725 267
rect 781 539 782 541
rect 784 539 785 541
rect 781 545 782 547
rect 784 545 785 547
rect 561 719 562 721
rect 564 719 565 721
rect 561 725 562 727
rect 564 725 565 727
rect 501 259 502 261
rect 504 259 505 261
rect 501 265 502 267
rect 504 265 505 267
rect 241 639 242 641
rect 244 639 245 641
rect 241 645 242 647
rect 244 645 245 647
rect 461 399 462 401
rect 464 399 465 401
rect 461 405 462 407
rect 464 405 465 407
rect 741 319 742 321
rect 744 319 745 321
rect 741 325 742 327
rect 744 325 745 327
rect 361 699 362 701
rect 364 699 365 701
rect 361 705 362 707
rect 364 705 365 707
rect 441 719 442 721
rect 444 719 445 721
rect 441 725 442 727
rect 444 725 445 727
rect 401 619 402 621
rect 404 619 405 621
rect 401 625 402 627
rect 404 625 405 627
rect 421 419 422 421
rect 424 419 425 421
rect 421 425 422 427
rect 424 425 425 427
rect 221 399 222 401
rect 224 399 225 401
rect 221 405 222 407
rect 224 405 225 407
rect 741 579 742 581
rect 744 579 745 581
rect 741 585 742 587
rect 744 585 745 587
rect 461 259 462 261
rect 464 259 465 261
rect 461 265 462 267
rect 464 265 465 267
rect 741 519 742 521
rect 744 519 745 521
rect 741 525 742 527
rect 744 525 745 527
rect 461 779 462 781
rect 464 779 465 781
rect 461 785 462 787
rect 464 785 465 787
rect 101 559 102 561
rect 104 559 105 561
rect 101 565 102 567
rect 104 565 105 567
rect 481 719 482 721
rect 484 719 485 721
rect 481 725 482 727
rect 484 725 485 727
rect 581 679 582 681
rect 584 679 585 681
rect 581 685 582 687
rect 584 685 585 687
rect 541 759 542 761
rect 544 759 545 761
rect 541 765 542 767
rect 544 765 545 767
rect 421 279 422 281
rect 424 279 425 281
rect 421 285 422 287
rect 424 285 425 287
rect 681 239 682 241
rect 684 239 685 241
rect 681 245 682 247
rect 684 245 685 247
rect 161 499 162 501
rect 164 499 165 501
rect 161 505 162 507
rect 164 505 165 507
rect 641 519 642 521
rect 644 519 645 521
rect 641 525 642 527
rect 644 525 645 527
rect 861 479 862 481
rect 864 479 865 481
rect 861 485 862 487
rect 864 485 865 487
rect 681 719 682 721
rect 684 719 685 721
rect 681 725 682 727
rect 684 725 685 727
rect 461 179 462 181
rect 464 179 465 181
rect 461 185 462 187
rect 464 185 465 187
rect 561 859 562 861
rect 564 859 565 861
rect 561 865 562 867
rect 564 865 565 867
rect 241 359 242 361
rect 244 359 245 361
rect 241 365 242 367
rect 244 365 245 367
rect 701 279 702 281
rect 704 279 705 281
rect 701 285 702 287
rect 704 285 705 287
rect 261 699 262 701
rect 264 699 265 701
rect 261 705 262 707
rect 264 705 265 707
rect 141 439 142 441
rect 144 439 145 441
rect 141 445 142 447
rect 144 445 145 447
rect 241 539 242 541
rect 244 539 245 541
rect 241 545 242 547
rect 244 545 245 547
rect 841 619 842 621
rect 844 619 845 621
rect 841 625 842 627
rect 844 625 845 627
rect 781 339 782 341
rect 784 339 785 341
rect 781 345 782 347
rect 784 345 785 347
rect 221 419 222 421
rect 224 419 225 421
rect 221 425 222 427
rect 224 425 225 427
rect 561 279 562 281
rect 564 279 565 281
rect 561 285 562 287
rect 564 285 565 287
rect 461 419 462 421
rect 464 419 465 421
rect 461 425 462 427
rect 464 425 465 427
rect 421 699 422 701
rect 424 699 425 701
rect 421 705 422 707
rect 424 705 425 707
rect 141 559 142 561
rect 144 559 145 561
rect 141 565 142 567
rect 144 565 145 567
rect 681 499 682 501
rect 684 499 685 501
rect 681 505 682 507
rect 684 505 685 507
rect 821 559 822 561
rect 824 559 825 561
rect 821 565 822 567
rect 824 565 825 567
rect 561 319 562 321
rect 564 319 565 321
rect 561 325 562 327
rect 564 325 565 327
rect 841 579 842 581
rect 844 579 845 581
rect 841 585 842 587
rect 844 585 845 587
rect 561 759 562 761
rect 564 759 565 761
rect 561 765 562 767
rect 564 765 565 767
rect 701 679 702 681
rect 704 679 705 681
rect 701 685 702 687
rect 704 685 705 687
rect 441 599 442 601
rect 444 599 445 601
rect 441 605 442 607
rect 444 605 445 607
rect 501 779 502 781
rect 504 779 505 781
rect 501 785 502 787
rect 504 785 505 787
rect 501 219 502 221
rect 504 219 505 221
rect 501 225 502 227
rect 504 225 505 227
rect 261 459 262 461
rect 264 459 265 461
rect 261 465 262 467
rect 264 465 265 467
rect 541 259 542 261
rect 544 259 545 261
rect 541 265 542 267
rect 544 265 545 267
rect 661 279 662 281
rect 664 279 665 281
rect 661 285 662 287
rect 664 285 665 287
rect 621 219 622 221
rect 624 219 625 221
rect 621 225 622 227
rect 624 225 625 227
rect 721 279 722 281
rect 724 279 725 281
rect 721 285 722 287
rect 724 285 725 287
rect 681 559 682 561
rect 684 559 685 561
rect 681 565 682 567
rect 684 565 685 567
rect 701 619 702 621
rect 704 619 705 621
rect 701 625 702 627
rect 704 625 705 627
rect 821 779 822 781
rect 824 779 825 781
rect 821 785 822 787
rect 824 785 825 787
rect 241 419 242 421
rect 244 419 245 421
rect 241 425 242 427
rect 244 425 245 427
rect 341 299 342 301
rect 344 299 345 301
rect 341 305 342 307
rect 344 305 345 307
rect 581 159 582 161
rect 584 159 585 161
rect 581 165 582 167
rect 584 165 585 167
rect 501 679 502 681
rect 504 679 505 681
rect 501 685 502 687
rect 504 685 505 687
rect 821 399 822 401
rect 824 399 825 401
rect 821 405 822 407
rect 824 405 825 407
rect 421 499 422 501
rect 424 499 425 501
rect 421 505 422 507
rect 424 505 425 507
rect 701 419 702 421
rect 704 419 705 421
rect 701 425 702 427
rect 704 425 705 427
rect 621 199 622 201
rect 624 199 625 201
rect 621 205 622 207
rect 624 205 625 207
rect 481 219 482 221
rect 484 219 485 221
rect 481 225 482 227
rect 484 225 485 227
rect 141 539 142 541
rect 144 539 145 541
rect 141 545 142 547
rect 144 545 145 547
rect 241 659 242 661
rect 244 659 245 661
rect 241 665 242 667
rect 244 665 245 667
rect 541 199 542 201
rect 544 199 545 201
rect 541 205 542 207
rect 544 205 545 207
rect 381 419 382 421
rect 384 419 385 421
rect 381 425 382 427
rect 384 425 385 427
rect 441 819 442 821
rect 444 819 445 821
rect 441 825 442 827
rect 444 825 445 827
rect 281 399 282 401
rect 284 399 285 401
rect 281 405 282 407
rect 284 405 285 407
rect 661 239 662 241
rect 664 239 665 241
rect 661 245 662 247
rect 664 245 665 247
rect 221 599 222 601
rect 224 599 225 601
rect 221 605 222 607
rect 224 605 225 607
rect 461 299 462 301
rect 464 299 465 301
rect 461 305 462 307
rect 464 305 465 307
rect 181 419 182 421
rect 184 419 185 421
rect 181 425 182 427
rect 184 425 185 427
rect 381 259 382 261
rect 384 259 385 261
rect 381 265 382 267
rect 384 265 385 267
rect 301 319 302 321
rect 304 319 305 321
rect 301 325 302 327
rect 304 325 305 327
rect 181 559 182 561
rect 184 559 185 561
rect 181 565 182 567
rect 184 565 185 567
rect 381 679 382 681
rect 384 679 385 681
rect 381 685 382 687
rect 384 685 385 687
rect 841 499 842 501
rect 844 499 845 501
rect 841 505 842 507
rect 844 505 845 507
rect 461 639 462 641
rect 464 639 465 641
rect 461 645 462 647
rect 464 645 465 647
rect 521 639 522 641
rect 524 639 525 641
rect 521 645 522 647
rect 524 645 525 647
rect 761 359 762 361
rect 764 359 765 361
rect 761 365 762 367
rect 764 365 765 367
rect 341 779 342 781
rect 344 779 345 781
rect 341 785 342 787
rect 344 785 345 787
rect 621 439 622 441
rect 624 439 625 441
rect 621 445 622 447
rect 624 445 625 447
rect 521 279 522 281
rect 524 279 525 281
rect 521 285 522 287
rect 524 285 525 287
rect 501 399 502 401
rect 504 399 505 401
rect 501 405 502 407
rect 504 405 505 407
rect 341 579 342 581
rect 344 579 345 581
rect 341 585 342 587
rect 344 585 345 587
rect 821 479 822 481
rect 824 479 825 481
rect 821 485 822 487
rect 824 485 825 487
rect 541 479 542 481
rect 544 479 545 481
rect 541 485 542 487
rect 544 485 545 487
rect 341 379 342 381
rect 344 379 345 381
rect 341 385 342 387
rect 344 385 345 387
rect 461 459 462 461
rect 464 459 465 461
rect 461 465 462 467
rect 464 465 465 467
rect 561 239 562 241
rect 564 239 565 241
rect 561 245 562 247
rect 564 245 565 247
rect 601 779 602 781
rect 604 779 605 781
rect 601 785 602 787
rect 604 785 605 787
rect 501 659 502 661
rect 504 659 505 661
rect 501 665 502 667
rect 504 665 505 667
rect 281 479 282 481
rect 284 479 285 481
rect 281 485 282 487
rect 284 485 285 487
rect 781 439 782 441
rect 784 439 785 441
rect 781 445 782 447
rect 784 445 785 447
rect 481 239 482 241
rect 484 239 485 241
rect 481 245 482 247
rect 484 245 485 247
rect 701 739 702 741
rect 704 739 705 741
rect 701 745 702 747
rect 704 745 705 747
rect 541 399 542 401
rect 544 399 545 401
rect 541 405 542 407
rect 544 405 545 407
rect 441 159 442 161
rect 444 159 445 161
rect 441 165 442 167
rect 444 165 445 167
rect 121 599 122 601
rect 124 599 125 601
rect 121 605 122 607
rect 124 605 125 607
rect 701 579 702 581
rect 704 579 705 581
rect 701 585 702 587
rect 704 585 705 587
rect 461 539 462 541
rect 464 539 465 541
rect 461 545 462 547
rect 464 545 465 547
rect 401 299 402 301
rect 404 299 405 301
rect 401 305 402 307
rect 404 305 405 307
rect 321 319 322 321
rect 324 319 325 321
rect 321 325 322 327
rect 324 325 325 327
rect 261 579 262 581
rect 264 579 265 581
rect 261 585 262 587
rect 264 585 265 587
rect 561 599 562 601
rect 564 599 565 601
rect 561 605 562 607
rect 564 605 565 607
rect 641 179 642 181
rect 644 179 645 181
rect 641 185 642 187
rect 644 185 645 187
rect 721 759 722 761
rect 724 759 725 761
rect 721 765 722 767
rect 724 765 725 767
rect 121 459 122 461
rect 124 459 125 461
rect 121 465 122 467
rect 124 465 125 467
rect 401 599 402 601
rect 404 599 405 601
rect 401 605 402 607
rect 404 605 405 607
rect 521 399 522 401
rect 524 399 525 401
rect 521 405 522 407
rect 524 405 525 407
rect 681 199 682 201
rect 684 199 685 201
rect 681 205 682 207
rect 684 205 685 207
rect 621 519 622 521
rect 624 519 625 521
rect 621 525 622 527
rect 624 525 625 527
rect 261 599 262 601
rect 264 599 265 601
rect 261 605 262 607
rect 264 605 265 607
rect 521 739 522 741
rect 524 739 525 741
rect 521 745 522 747
rect 524 745 525 747
rect 621 419 622 421
rect 624 419 625 421
rect 621 425 622 427
rect 624 425 625 427
rect 281 679 282 681
rect 284 679 285 681
rect 281 685 282 687
rect 284 685 285 687
rect 421 639 422 641
rect 424 639 425 641
rect 421 645 422 647
rect 424 645 425 647
rect 561 299 562 301
rect 564 299 565 301
rect 561 305 562 307
rect 564 305 565 307
rect 321 679 322 681
rect 324 679 325 681
rect 321 685 322 687
rect 324 685 325 687
rect 561 499 562 501
rect 564 499 565 501
rect 561 505 562 507
rect 564 505 565 507
rect 241 479 242 481
rect 244 479 245 481
rect 241 485 242 487
rect 244 485 245 487
rect 701 599 702 601
rect 704 599 705 601
rect 701 605 702 607
rect 704 605 705 607
rect 281 639 282 641
rect 284 639 285 641
rect 281 645 282 647
rect 284 645 285 647
rect 301 559 302 561
rect 304 559 305 561
rect 301 565 302 567
rect 304 565 305 567
rect 441 439 442 441
rect 444 439 445 441
rect 441 445 442 447
rect 444 445 445 447
rect 601 439 602 441
rect 604 439 605 441
rect 601 445 602 447
rect 604 445 605 447
rect 621 459 622 461
rect 624 459 625 461
rect 621 465 622 467
rect 624 465 625 467
rect 661 579 662 581
rect 664 579 665 581
rect 661 585 662 587
rect 664 585 665 587
rect 401 639 402 641
rect 404 639 405 641
rect 401 645 402 647
rect 404 645 405 647
rect 261 439 262 441
rect 264 439 265 441
rect 261 445 262 447
rect 264 445 265 447
rect 861 579 862 581
rect 864 579 865 581
rect 861 585 862 587
rect 864 585 865 587
rect 721 639 722 641
rect 724 639 725 641
rect 721 645 722 647
rect 724 645 725 647
rect 381 299 382 301
rect 384 299 385 301
rect 381 305 382 307
rect 384 305 385 307
rect 421 719 422 721
rect 424 719 425 721
rect 421 725 422 727
rect 424 725 425 727
rect 301 679 302 681
rect 304 679 305 681
rect 301 685 302 687
rect 304 685 305 687
rect 621 659 622 661
rect 624 659 625 661
rect 621 665 622 667
rect 624 665 625 667
rect 701 519 702 521
rect 704 519 705 521
rect 701 525 702 527
rect 704 525 705 527
rect 321 759 322 761
rect 324 759 325 761
rect 321 765 322 767
rect 324 765 325 767
rect 481 779 482 781
rect 484 779 485 781
rect 481 785 482 787
rect 484 785 485 787
rect 701 639 702 641
rect 704 639 705 641
rect 701 645 702 647
rect 704 645 705 647
rect 581 519 582 521
rect 584 519 585 521
rect 581 525 582 527
rect 584 525 585 527
rect 601 519 602 521
rect 604 519 605 521
rect 601 525 602 527
rect 604 525 605 527
rect 461 479 462 481
rect 464 479 465 481
rect 461 485 462 487
rect 464 485 465 487
rect 601 679 602 681
rect 604 679 605 681
rect 601 685 602 687
rect 604 685 605 687
rect 481 699 482 701
rect 484 699 485 701
rect 481 705 482 707
rect 484 705 485 707
rect 761 639 762 641
rect 764 639 765 641
rect 761 645 762 647
rect 764 645 765 647
rect 421 739 422 741
rect 424 739 425 741
rect 421 745 422 747
rect 424 745 425 747
rect 701 259 702 261
rect 704 259 705 261
rect 701 265 702 267
rect 704 265 705 267
rect 441 739 442 741
rect 444 739 445 741
rect 441 745 442 747
rect 444 745 445 747
rect 381 359 382 361
rect 384 359 385 361
rect 381 365 382 367
rect 384 365 385 367
rect 341 599 342 601
rect 344 599 345 601
rect 341 605 342 607
rect 344 605 345 607
rect 561 619 562 621
rect 564 619 565 621
rect 561 625 562 627
rect 564 625 565 627
rect 641 439 642 441
rect 644 439 645 441
rect 641 445 642 447
rect 644 445 645 447
rect 321 279 322 281
rect 324 279 325 281
rect 321 285 322 287
rect 324 285 325 287
rect 661 359 662 361
rect 664 359 665 361
rect 661 365 662 367
rect 664 365 665 367
rect 301 539 302 541
rect 304 539 305 541
rect 301 545 302 547
rect 304 545 305 547
rect 401 699 402 701
rect 404 699 405 701
rect 401 705 402 707
rect 404 705 405 707
rect 621 479 622 481
rect 624 479 625 481
rect 621 485 622 487
rect 624 485 625 487
rect 541 219 542 221
rect 544 219 545 221
rect 541 225 542 227
rect 544 225 545 227
rect 581 339 582 341
rect 584 339 585 341
rect 581 345 582 347
rect 584 345 585 347
rect 501 699 502 701
rect 504 699 505 701
rect 501 705 502 707
rect 504 705 505 707
rect 481 439 482 441
rect 484 439 485 441
rect 481 445 482 447
rect 484 445 485 447
rect 721 539 722 541
rect 724 539 725 541
rect 721 545 722 547
rect 724 545 725 547
rect 301 619 302 621
rect 304 619 305 621
rect 301 625 302 627
rect 304 625 305 627
rect 861 599 862 601
rect 864 599 865 601
rect 861 605 862 607
rect 864 605 865 607
rect 521 679 522 681
rect 524 679 525 681
rect 521 685 522 687
rect 524 685 525 687
rect 761 539 762 541
rect 764 539 765 541
rect 761 545 762 547
rect 764 545 765 547
rect 221 639 222 641
rect 224 639 225 641
rect 221 645 222 647
rect 224 645 225 647
rect 301 499 302 501
rect 304 499 305 501
rect 301 505 302 507
rect 304 505 305 507
rect 401 279 402 281
rect 404 279 405 281
rect 401 285 402 287
rect 404 285 405 287
rect 441 659 442 661
rect 444 659 445 661
rect 441 665 442 667
rect 444 665 445 667
rect 541 599 542 601
rect 544 599 545 601
rect 541 605 542 607
rect 544 605 545 607
rect 361 539 362 541
rect 364 539 365 541
rect 361 545 362 547
rect 364 545 365 547
rect 341 799 342 801
rect 344 799 345 801
rect 341 805 342 807
rect 344 805 345 807
rect 581 639 582 641
rect 584 639 585 641
rect 581 645 582 647
rect 584 645 585 647
rect 501 339 502 341
rect 504 339 505 341
rect 501 345 502 347
rect 504 345 505 347
rect 201 639 202 641
rect 204 639 205 641
rect 201 645 202 647
rect 204 645 205 647
rect 661 799 662 801
rect 664 799 665 801
rect 661 805 662 807
rect 664 805 665 807
rect 161 479 162 481
rect 164 479 165 481
rect 161 485 162 487
rect 164 485 165 487
rect 301 359 302 361
rect 304 359 305 361
rect 301 365 302 367
rect 304 365 305 367
rect 421 539 422 541
rect 424 539 425 541
rect 421 545 422 547
rect 424 545 425 547
rect 621 539 622 541
rect 624 539 625 541
rect 621 545 622 547
rect 624 545 625 547
rect 461 319 462 321
rect 464 319 465 321
rect 461 325 462 327
rect 464 325 465 327
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect 521 299 522 301
rect 524 299 525 301
rect 521 305 522 307
rect 524 305 525 307
rect 641 359 642 361
rect 644 359 645 361
rect 641 365 642 367
rect 644 365 645 367
rect 221 539 222 541
rect 224 539 225 541
rect 221 545 222 547
rect 224 545 225 547
rect 401 459 402 461
rect 404 459 405 461
rect 401 465 402 467
rect 404 465 405 467
rect 641 599 642 601
rect 644 599 645 601
rect 641 605 642 607
rect 644 605 645 607
rect 881 559 882 561
rect 884 559 885 561
rect 881 565 882 567
rect 884 565 885 567
rect 341 339 342 341
rect 344 339 345 341
rect 341 345 342 347
rect 344 345 345 347
rect 701 439 702 441
rect 704 439 705 441
rect 701 445 702 447
rect 704 445 705 447
rect 421 779 422 781
rect 424 779 425 781
rect 421 785 422 787
rect 424 785 425 787
rect 361 299 362 301
rect 364 299 365 301
rect 361 305 362 307
rect 364 305 365 307
rect 541 619 542 621
rect 544 619 545 621
rect 541 625 542 627
rect 544 625 545 627
rect 361 399 362 401
rect 364 399 365 401
rect 361 405 362 407
rect 364 405 365 407
rect 261 619 262 621
rect 264 619 265 621
rect 261 625 262 627
rect 264 625 265 627
rect 641 479 642 481
rect 644 479 645 481
rect 641 485 642 487
rect 644 485 645 487
rect 641 639 642 641
rect 644 639 645 641
rect 641 645 642 647
rect 644 645 645 647
rect 401 499 402 501
rect 404 499 405 501
rect 401 505 402 507
rect 404 505 405 507
rect 581 739 582 741
rect 584 739 585 741
rect 581 745 582 747
rect 584 745 585 747
rect 141 479 142 481
rect 144 479 145 481
rect 141 485 142 487
rect 144 485 145 487
rect 661 739 662 741
rect 664 739 665 741
rect 661 745 662 747
rect 664 745 665 747
rect 401 839 402 841
rect 404 839 405 841
rect 401 845 402 847
rect 404 845 405 847
rect 381 219 382 221
rect 384 219 385 221
rect 381 225 382 227
rect 384 225 385 227
rect 341 639 342 641
rect 344 639 345 641
rect 341 645 342 647
rect 344 645 345 647
rect 201 419 202 421
rect 204 419 205 421
rect 201 425 202 427
rect 204 425 205 427
rect 761 559 762 561
rect 764 559 765 561
rect 761 565 762 567
rect 764 565 765 567
rect 301 279 302 281
rect 304 279 305 281
rect 301 285 302 287
rect 304 285 305 287
rect 181 619 182 621
rect 184 619 185 621
rect 181 625 182 627
rect 184 625 185 627
rect 421 519 422 521
rect 424 519 425 521
rect 421 525 422 527
rect 424 525 425 527
rect 541 339 542 341
rect 544 339 545 341
rect 541 345 542 347
rect 544 345 545 347
rect 641 379 642 381
rect 644 379 645 381
rect 641 385 642 387
rect 644 385 645 387
rect 801 579 802 581
rect 804 579 805 581
rect 801 585 802 587
rect 804 585 805 587
rect 241 599 242 601
rect 244 599 245 601
rect 241 605 242 607
rect 244 605 245 607
rect 121 559 122 561
rect 124 559 125 561
rect 121 565 122 567
rect 124 565 125 567
rect 801 479 802 481
rect 804 479 805 481
rect 801 485 802 487
rect 804 485 805 487
rect 621 579 622 581
rect 624 579 625 581
rect 621 585 622 587
rect 624 585 625 587
rect 781 559 782 561
rect 784 559 785 561
rect 781 565 782 567
rect 784 565 785 567
rect 841 479 842 481
rect 844 479 845 481
rect 841 485 842 487
rect 844 485 845 487
rect 601 479 602 481
rect 604 479 605 481
rect 601 485 602 487
rect 604 485 605 487
rect 521 799 522 801
rect 524 799 525 801
rect 521 805 522 807
rect 524 805 525 807
rect 481 199 482 201
rect 484 199 485 201
rect 481 205 482 207
rect 484 205 485 207
rect 561 199 562 201
rect 564 199 565 201
rect 561 205 562 207
rect 564 205 565 207
rect 721 399 722 401
rect 724 399 725 401
rect 721 405 722 407
rect 724 405 725 407
rect 281 419 282 421
rect 284 419 285 421
rect 281 425 282 427
rect 284 425 285 427
rect 821 419 822 421
rect 824 419 825 421
rect 821 425 822 427
rect 824 425 825 427
rect 601 239 602 241
rect 604 239 605 241
rect 601 245 602 247
rect 604 245 605 247
rect 621 339 622 341
rect 624 339 625 341
rect 621 345 622 347
rect 624 345 625 347
rect 581 179 582 181
rect 584 179 585 181
rect 581 185 582 187
rect 584 185 585 187
rect 721 619 722 621
rect 724 619 725 621
rect 721 625 722 627
rect 724 625 725 627
rect 461 359 462 361
rect 464 359 465 361
rect 461 365 462 367
rect 464 365 465 367
rect 461 379 462 381
rect 464 379 465 381
rect 461 385 462 387
rect 464 385 465 387
rect 781 399 782 401
rect 784 399 785 401
rect 781 405 782 407
rect 784 405 785 407
rect 601 579 602 581
rect 604 579 605 581
rect 601 585 602 587
rect 604 585 605 587
rect 761 339 762 341
rect 764 339 765 341
rect 761 345 762 347
rect 764 345 765 347
rect 621 599 622 601
rect 624 599 625 601
rect 621 605 622 607
rect 624 605 625 607
rect 561 819 562 821
rect 564 819 565 821
rect 561 825 562 827
rect 564 825 565 827
rect 481 679 482 681
rect 484 679 485 681
rect 481 685 482 687
rect 484 685 485 687
rect 341 519 342 521
rect 344 519 345 521
rect 341 525 342 527
rect 344 525 345 527
rect 181 439 182 441
rect 184 439 185 441
rect 181 445 182 447
rect 184 445 185 447
rect 781 579 782 581
rect 784 579 785 581
rect 781 585 782 587
rect 784 585 785 587
rect 641 679 642 681
rect 644 679 645 681
rect 641 685 642 687
rect 644 685 645 687
rect 701 319 702 321
rect 704 319 705 321
rect 701 325 702 327
rect 704 325 705 327
rect 341 419 342 421
rect 344 419 345 421
rect 341 425 342 427
rect 344 425 345 427
rect 841 599 842 601
rect 844 599 845 601
rect 841 605 842 607
rect 844 605 845 607
rect 301 639 302 641
rect 304 639 305 641
rect 301 645 302 647
rect 304 645 305 647
rect 501 639 502 641
rect 504 639 505 641
rect 501 645 502 647
rect 504 645 505 647
rect 441 519 442 521
rect 444 519 445 521
rect 441 525 442 527
rect 444 525 445 527
rect 321 559 322 561
rect 324 559 325 561
rect 321 565 322 567
rect 324 565 325 567
rect 481 379 482 381
rect 484 379 485 381
rect 481 385 482 387
rect 484 385 485 387
rect 701 479 702 481
rect 704 479 705 481
rect 701 485 702 487
rect 704 485 705 487
rect 381 439 382 441
rect 384 439 385 441
rect 381 445 382 447
rect 384 445 385 447
rect 461 239 462 241
rect 464 239 465 241
rect 461 245 462 247
rect 464 245 465 247
rect 401 359 402 361
rect 404 359 405 361
rect 401 365 402 367
rect 404 365 405 367
rect 601 719 602 721
rect 604 719 605 721
rect 601 725 602 727
rect 604 725 605 727
rect 461 699 462 701
rect 464 699 465 701
rect 461 705 462 707
rect 464 705 465 707
rect 481 559 482 561
rect 484 559 485 561
rect 481 565 482 567
rect 484 565 485 567
rect 661 759 662 761
rect 664 759 665 761
rect 661 765 662 767
rect 664 765 665 767
rect 381 739 382 741
rect 384 739 385 741
rect 381 745 382 747
rect 384 745 385 747
rect 681 759 682 761
rect 684 759 685 761
rect 681 765 682 767
rect 684 765 685 767
rect 641 239 642 241
rect 644 239 645 241
rect 641 245 642 247
rect 644 245 645 247
rect 741 499 742 501
rect 744 499 745 501
rect 741 505 742 507
rect 744 505 745 507
rect 381 699 382 701
rect 384 699 385 701
rect 381 705 382 707
rect 384 705 385 707
rect 381 579 382 581
rect 384 579 385 581
rect 381 585 382 587
rect 384 585 385 587
rect 721 339 722 341
rect 724 339 725 341
rect 721 345 722 347
rect 724 345 725 347
rect 401 179 402 181
rect 404 179 405 181
rect 401 185 402 187
rect 404 185 405 187
rect 381 559 382 561
rect 384 559 385 561
rect 381 565 382 567
rect 384 565 385 567
rect 521 319 522 321
rect 524 319 525 321
rect 521 325 522 327
rect 524 325 525 327
rect 681 299 682 301
rect 684 299 685 301
rect 681 305 682 307
rect 684 305 685 307
rect 661 259 662 261
rect 664 259 665 261
rect 661 265 662 267
rect 664 265 665 267
rect 461 199 462 201
rect 464 199 465 201
rect 461 205 462 207
rect 464 205 465 207
rect 221 619 222 621
rect 224 619 225 621
rect 221 625 222 627
rect 224 625 225 627
rect 381 819 382 821
rect 384 819 385 821
rect 381 825 382 827
rect 384 825 385 827
rect 621 639 622 641
rect 624 639 625 641
rect 621 645 622 647
rect 624 645 625 647
rect 421 439 422 441
rect 424 439 425 441
rect 421 445 422 447
rect 424 445 425 447
rect 321 519 322 521
rect 324 519 325 521
rect 321 525 322 527
rect 324 525 325 527
rect 401 579 402 581
rect 404 579 405 581
rect 401 585 402 587
rect 404 585 405 587
rect 381 799 382 801
rect 384 799 385 801
rect 381 805 382 807
rect 384 805 385 807
rect 601 599 602 601
rect 604 599 605 601
rect 601 605 602 607
rect 604 605 605 607
rect 541 739 542 741
rect 544 739 545 741
rect 541 745 542 747
rect 544 745 545 747
rect 481 619 482 621
rect 484 619 485 621
rect 481 625 482 627
rect 484 625 485 627
rect 801 519 802 521
rect 804 519 805 521
rect 801 525 802 527
rect 804 525 805 527
rect 561 679 562 681
rect 564 679 565 681
rect 561 685 562 687
rect 564 685 565 687
rect 581 619 582 621
rect 584 619 585 621
rect 581 625 582 627
rect 584 625 585 627
rect 241 399 242 401
rect 244 399 245 401
rect 241 405 242 407
rect 244 405 245 407
rect 601 359 602 361
rect 604 359 605 361
rect 601 365 602 367
rect 604 365 605 367
rect 521 879 522 881
rect 524 879 525 881
rect 521 885 522 887
rect 524 885 525 887
rect 541 379 542 381
rect 544 379 545 381
rect 541 385 542 387
rect 544 385 545 387
rect 221 579 222 581
rect 224 579 225 581
rect 221 585 222 587
rect 224 585 225 587
rect 681 739 682 741
rect 684 739 685 741
rect 681 745 682 747
rect 684 745 685 747
rect 401 479 402 481
rect 404 479 405 481
rect 401 485 402 487
rect 404 485 405 487
rect 761 619 762 621
rect 764 619 765 621
rect 761 625 762 627
rect 764 625 765 627
rect 601 759 602 761
rect 604 759 605 761
rect 601 765 602 767
rect 604 765 605 767
rect 601 659 602 661
rect 604 659 605 661
rect 601 665 602 667
rect 604 665 605 667
rect 461 759 462 761
rect 464 759 465 761
rect 461 765 462 767
rect 464 765 465 767
rect 601 319 602 321
rect 604 319 605 321
rect 601 325 602 327
rect 604 325 605 327
rect 701 379 702 381
rect 704 379 705 381
rect 701 385 702 387
rect 704 385 705 387
rect 701 719 702 721
rect 704 719 705 721
rect 701 725 702 727
rect 704 725 705 727
rect 681 779 682 781
rect 684 779 685 781
rect 681 785 682 787
rect 684 785 685 787
rect 541 719 542 721
rect 544 719 545 721
rect 541 725 542 727
rect 544 725 545 727
rect 281 659 282 661
rect 284 659 285 661
rect 281 665 282 667
rect 284 665 285 667
rect 761 439 762 441
rect 764 439 765 441
rect 761 445 762 447
rect 764 445 765 447
rect 501 499 502 501
rect 504 499 505 501
rect 501 505 502 507
rect 504 505 505 507
rect 241 459 242 461
rect 244 459 245 461
rect 241 465 242 467
rect 244 465 245 467
rect 321 399 322 401
rect 324 399 325 401
rect 321 405 322 407
rect 324 405 325 407
rect 541 859 542 861
rect 544 859 545 861
rect 541 865 542 867
rect 544 865 545 867
rect 261 419 262 421
rect 264 419 265 421
rect 261 425 262 427
rect 264 425 265 427
rect 681 619 682 621
rect 684 619 685 621
rect 681 625 682 627
rect 684 625 685 627
rect 321 299 322 301
rect 324 299 325 301
rect 321 305 322 307
rect 324 305 325 307
rect 641 659 642 661
rect 644 659 645 661
rect 641 665 642 667
rect 644 665 645 667
rect 661 719 662 721
rect 664 719 665 721
rect 661 725 662 727
rect 664 725 665 727
rect 581 499 582 501
rect 584 499 585 501
rect 581 505 582 507
rect 584 505 585 507
rect 441 479 442 481
rect 444 479 445 481
rect 441 485 442 487
rect 444 485 445 487
rect 681 799 682 801
rect 684 799 685 801
rect 681 805 682 807
rect 684 805 685 807
rect 621 359 622 361
rect 624 359 625 361
rect 621 365 622 367
rect 624 365 625 367
rect 501 479 502 481
rect 504 479 505 481
rect 501 485 502 487
rect 504 485 505 487
rect 281 699 282 701
rect 284 699 285 701
rect 281 705 282 707
rect 284 705 285 707
rect 201 599 202 601
rect 204 599 205 601
rect 201 605 202 607
rect 204 605 205 607
rect 761 679 762 681
rect 764 679 765 681
rect 761 685 762 687
rect 764 685 765 687
rect 581 539 582 541
rect 584 539 585 541
rect 581 545 582 547
rect 584 545 585 547
rect 121 539 122 541
rect 124 539 125 541
rect 121 545 122 547
rect 124 545 125 547
rect 181 599 182 601
rect 184 599 185 601
rect 181 605 182 607
rect 184 605 185 607
rect 521 379 522 381
rect 524 379 525 381
rect 521 385 522 387
rect 524 385 525 387
rect 501 439 502 441
rect 504 439 505 441
rect 501 445 502 447
rect 504 445 505 447
rect 341 279 342 281
rect 344 279 345 281
rect 341 285 342 287
rect 344 285 345 287
rect 441 419 442 421
rect 444 419 445 421
rect 441 425 442 427
rect 444 425 445 427
rect 741 539 742 541
rect 744 539 745 541
rect 741 545 742 547
rect 744 545 745 547
rect 541 879 542 881
rect 544 879 545 881
rect 541 885 542 887
rect 544 885 545 887
rect 461 279 462 281
rect 464 279 465 281
rect 461 285 462 287
rect 464 285 465 287
rect 381 539 382 541
rect 384 539 385 541
rect 381 545 382 547
rect 384 545 385 547
rect 681 539 682 541
rect 684 539 685 541
rect 681 545 682 547
rect 684 545 685 547
rect 501 299 502 301
rect 504 299 505 301
rect 501 305 502 307
rect 504 305 505 307
rect 361 319 362 321
rect 364 319 365 321
rect 361 325 362 327
rect 364 325 365 327
rect 521 339 522 341
rect 524 339 525 341
rect 521 345 522 347
rect 524 345 525 347
rect 681 319 682 321
rect 684 319 685 321
rect 681 325 682 327
rect 684 325 685 327
rect 541 699 542 701
rect 544 699 545 701
rect 541 705 542 707
rect 544 705 545 707
rect 421 619 422 621
rect 424 619 425 621
rect 421 625 422 627
rect 424 625 425 627
rect 661 559 662 561
rect 664 559 665 561
rect 661 565 662 567
rect 664 565 665 567
rect 541 299 542 301
rect 544 299 545 301
rect 541 305 542 307
rect 544 305 545 307
rect 541 799 542 801
rect 544 799 545 801
rect 541 805 542 807
rect 544 805 545 807
rect 301 459 302 461
rect 304 459 305 461
rect 301 465 302 467
rect 304 465 305 467
rect 581 599 582 601
rect 584 599 585 601
rect 581 605 582 607
rect 584 605 585 607
rect 381 779 382 781
rect 384 779 385 781
rect 381 785 382 787
rect 384 785 385 787
rect 481 479 482 481
rect 484 479 485 481
rect 481 485 482 487
rect 484 485 485 487
rect 401 399 402 401
rect 404 399 405 401
rect 401 405 402 407
rect 404 405 405 407
rect 581 299 582 301
rect 584 299 585 301
rect 581 305 582 307
rect 584 305 585 307
rect 661 419 662 421
rect 664 419 665 421
rect 661 425 662 427
rect 664 425 665 427
rect 201 399 202 401
rect 204 399 205 401
rect 201 405 202 407
rect 204 405 205 407
rect 521 239 522 241
rect 524 239 525 241
rect 521 245 522 247
rect 524 245 525 247
rect 341 659 342 661
rect 344 659 345 661
rect 341 665 342 667
rect 344 665 345 667
rect 801 659 802 661
rect 804 659 805 661
rect 801 665 802 667
rect 804 665 805 667
rect 301 519 302 521
rect 304 519 305 521
rect 301 525 302 527
rect 304 525 305 527
rect 661 299 662 301
rect 664 299 665 301
rect 661 305 662 307
rect 664 305 665 307
rect 601 499 602 501
rect 604 499 605 501
rect 601 505 602 507
rect 604 505 605 507
rect 341 239 342 241
rect 344 239 345 241
rect 341 245 342 247
rect 344 245 345 247
rect 741 419 742 421
rect 744 419 745 421
rect 741 425 742 427
rect 744 425 745 427
rect 581 859 582 861
rect 584 859 585 861
rect 581 865 582 867
rect 584 865 585 867
rect 201 459 202 461
rect 204 459 205 461
rect 201 465 202 467
rect 204 465 205 467
rect 721 379 722 381
rect 724 379 725 381
rect 721 385 722 387
rect 724 385 725 387
rect 421 759 422 761
rect 424 759 425 761
rect 421 765 422 767
rect 424 765 425 767
rect 641 759 642 761
rect 644 759 645 761
rect 641 765 642 767
rect 644 765 645 767
rect 581 379 582 381
rect 584 379 585 381
rect 581 385 582 387
rect 584 385 585 387
rect 561 839 562 841
rect 564 839 565 841
rect 561 845 562 847
rect 564 845 565 847
rect 381 619 382 621
rect 384 619 385 621
rect 381 625 382 627
rect 384 625 385 627
rect 681 459 682 461
rect 684 459 685 461
rect 681 465 682 467
rect 684 465 685 467
rect 461 559 462 561
rect 464 559 465 561
rect 461 565 462 567
rect 464 565 465 567
rect 621 319 622 321
rect 624 319 625 321
rect 621 325 622 327
rect 624 325 625 327
rect 501 359 502 361
rect 504 359 505 361
rect 501 365 502 367
rect 504 365 505 367
rect 601 299 602 301
rect 604 299 605 301
rect 601 305 602 307
rect 604 305 605 307
rect 441 399 442 401
rect 444 399 445 401
rect 441 405 442 407
rect 444 405 445 407
rect 401 719 402 721
rect 404 719 405 721
rect 401 725 402 727
rect 404 725 405 727
rect 881 579 882 581
rect 884 579 885 581
rect 881 585 882 587
rect 884 585 885 587
rect 321 739 322 741
rect 324 739 325 741
rect 321 745 322 747
rect 324 745 325 747
rect 581 839 582 841
rect 584 839 585 841
rect 581 845 582 847
rect 584 845 585 847
rect 521 479 522 481
rect 524 479 525 481
rect 521 485 522 487
rect 524 485 525 487
rect 301 759 302 761
rect 304 759 305 761
rect 301 765 302 767
rect 304 765 305 767
rect 841 519 842 521
rect 844 519 845 521
rect 841 525 842 527
rect 844 525 845 527
rect 401 199 402 201
rect 404 199 405 201
rect 401 205 402 207
rect 404 205 405 207
rect 561 379 562 381
rect 564 379 565 381
rect 561 385 562 387
rect 564 385 565 387
rect 361 239 362 241
rect 364 239 365 241
rect 361 245 362 247
rect 364 245 365 247
rect 381 499 382 501
rect 384 499 385 501
rect 381 505 382 507
rect 384 505 385 507
rect 561 519 562 521
rect 564 519 565 521
rect 561 525 562 527
rect 564 525 565 527
rect 161 639 162 641
rect 164 639 165 641
rect 161 645 162 647
rect 164 645 165 647
rect 581 459 582 461
rect 584 459 585 461
rect 581 465 582 467
rect 584 465 585 467
rect 481 499 482 501
rect 484 499 485 501
rect 481 505 482 507
rect 484 505 485 507
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect 661 679 662 681
rect 664 679 665 681
rect 661 685 662 687
rect 664 685 665 687
rect 481 599 482 601
rect 484 599 485 601
rect 481 605 482 607
rect 484 605 485 607
rect 241 719 242 721
rect 244 719 245 721
rect 241 725 242 727
rect 244 725 245 727
rect 341 359 342 361
rect 344 359 345 361
rect 341 365 342 367
rect 344 365 345 367
rect 361 639 362 641
rect 364 639 365 641
rect 361 645 362 647
rect 364 645 365 647
rect 401 679 402 681
rect 404 679 405 681
rect 401 685 402 687
rect 404 685 405 687
rect 581 359 582 361
rect 584 359 585 361
rect 581 365 582 367
rect 584 365 585 367
rect 621 279 622 281
rect 624 279 625 281
rect 621 285 622 287
rect 624 285 625 287
rect 601 179 602 181
rect 604 179 605 181
rect 601 185 602 187
rect 604 185 605 187
rect 681 639 682 641
rect 684 639 685 641
rect 681 645 682 647
rect 684 645 685 647
rect 501 159 502 161
rect 504 159 505 161
rect 501 165 502 167
rect 504 165 505 167
rect 561 339 562 341
rect 564 339 565 341
rect 561 345 562 347
rect 564 345 565 347
rect 681 339 682 341
rect 684 339 685 341
rect 681 345 682 347
rect 684 345 685 347
rect 521 899 522 901
rect 524 899 525 901
rect 521 905 522 907
rect 524 905 525 907
rect 581 279 582 281
rect 584 279 585 281
rect 581 285 582 287
rect 584 285 585 287
rect 561 779 562 781
rect 564 779 565 781
rect 561 785 562 787
rect 564 785 565 787
rect 401 379 402 381
rect 404 379 405 381
rect 401 385 402 387
rect 404 385 405 387
rect 281 359 282 361
rect 284 359 285 361
rect 281 365 282 367
rect 284 365 285 367
rect 441 639 442 641
rect 444 639 445 641
rect 441 645 442 647
rect 444 645 445 647
rect 561 179 562 181
rect 564 179 565 181
rect 561 185 562 187
rect 564 185 565 187
rect 781 459 782 461
rect 784 459 785 461
rect 781 465 782 467
rect 784 465 785 467
rect 861 439 862 441
rect 864 439 865 441
rect 861 445 862 447
rect 864 445 865 447
rect 781 599 782 601
rect 784 599 785 601
rect 781 605 782 607
rect 784 605 785 607
rect 361 459 362 461
rect 364 459 365 461
rect 361 465 362 467
rect 364 465 365 467
rect 401 519 402 521
rect 404 519 405 521
rect 401 525 402 527
rect 404 525 405 527
rect 741 339 742 341
rect 744 339 745 341
rect 741 345 742 347
rect 744 345 745 347
rect 821 539 822 541
rect 824 539 825 541
rect 821 545 822 547
rect 824 545 825 547
rect 441 259 442 261
rect 444 259 445 261
rect 441 265 442 267
rect 444 265 445 267
rect 341 459 342 461
rect 344 459 345 461
rect 341 465 342 467
rect 344 465 345 467
rect 661 399 662 401
rect 664 399 665 401
rect 661 405 662 407
rect 664 405 665 407
rect 561 559 562 561
rect 564 559 565 561
rect 561 565 562 567
rect 564 565 565 567
rect 601 259 602 261
rect 604 259 605 261
rect 601 265 602 267
rect 604 265 605 267
rect 781 479 782 481
rect 784 479 785 481
rect 781 485 782 487
rect 784 485 785 487
rect 441 219 442 221
rect 444 219 445 221
rect 441 225 442 227
rect 444 225 445 227
rect 201 559 202 561
rect 204 559 205 561
rect 201 565 202 567
rect 204 565 205 567
rect 181 459 182 461
rect 184 459 185 461
rect 181 465 182 467
rect 184 465 185 467
rect 301 779 302 781
rect 304 779 305 781
rect 301 785 302 787
rect 304 785 305 787
rect 661 699 662 701
rect 664 699 665 701
rect 661 705 662 707
rect 664 705 665 707
rect 601 379 602 381
rect 604 379 605 381
rect 601 385 602 387
rect 604 385 605 387
rect 621 239 622 241
rect 624 239 625 241
rect 621 245 622 247
rect 624 245 625 247
rect 721 699 722 701
rect 724 699 725 701
rect 721 705 722 707
rect 724 705 725 707
rect 421 299 422 301
rect 424 299 425 301
rect 421 305 422 307
rect 424 305 425 307
rect 181 399 182 401
rect 184 399 185 401
rect 181 405 182 407
rect 184 405 185 407
rect 421 239 422 241
rect 424 239 425 241
rect 421 245 422 247
rect 424 245 425 247
rect 521 499 522 501
rect 524 499 525 501
rect 521 505 522 507
rect 524 505 525 507
rect 681 419 682 421
rect 684 419 685 421
rect 681 425 682 427
rect 684 425 685 427
rect 361 479 362 481
rect 364 479 365 481
rect 361 485 362 487
rect 364 485 365 487
rect 761 579 762 581
rect 764 579 765 581
rect 761 585 762 587
rect 764 585 765 587
rect 601 639 602 641
rect 604 639 605 641
rect 601 645 602 647
rect 604 645 605 647
rect 301 399 302 401
rect 304 399 305 401
rect 301 405 302 407
rect 304 405 305 407
rect 201 479 202 481
rect 204 479 205 481
rect 201 485 202 487
rect 204 485 205 487
rect 661 479 662 481
rect 664 479 665 481
rect 661 485 662 487
rect 664 485 665 487
rect 741 559 742 561
rect 744 559 745 561
rect 741 565 742 567
rect 744 565 745 567
rect 721 599 722 601
rect 724 599 725 601
rect 721 605 722 607
rect 724 605 725 607
rect 641 739 642 741
rect 644 739 645 741
rect 641 745 642 747
rect 644 745 645 747
rect 301 339 302 341
rect 304 339 305 341
rect 301 345 302 347
rect 304 345 305 347
rect 721 319 722 321
rect 724 319 725 321
rect 721 325 722 327
rect 724 325 725 327
rect 241 739 242 741
rect 244 739 245 741
rect 241 745 242 747
rect 244 745 245 747
rect 481 879 482 881
rect 484 879 485 881
rect 481 885 482 887
rect 484 885 485 887
rect 561 439 562 441
rect 564 439 565 441
rect 561 445 562 447
rect 564 445 565 447
rect 481 359 482 361
rect 484 359 485 361
rect 481 365 482 367
rect 484 365 485 367
rect 601 539 602 541
rect 604 539 605 541
rect 601 545 602 547
rect 604 545 605 547
rect 661 519 662 521
rect 664 519 665 521
rect 661 525 662 527
rect 664 525 665 527
rect 361 359 362 361
rect 364 359 365 361
rect 361 365 362 367
rect 364 365 365 367
rect 221 379 222 381
rect 224 379 225 381
rect 221 385 222 387
rect 224 385 225 387
rect 821 619 822 621
rect 824 619 825 621
rect 821 625 822 627
rect 824 625 825 627
rect 681 279 682 281
rect 684 279 685 281
rect 681 285 682 287
rect 684 285 685 287
rect 361 679 362 681
rect 364 679 365 681
rect 361 685 362 687
rect 364 685 365 687
rect 361 659 362 661
rect 364 659 365 661
rect 361 665 362 667
rect 364 665 365 667
rect 161 459 162 461
rect 164 459 165 461
rect 161 465 162 467
rect 164 465 165 467
rect 481 519 482 521
rect 484 519 485 521
rect 481 525 482 527
rect 484 525 485 527
rect 361 499 362 501
rect 364 499 365 501
rect 361 505 362 507
rect 364 505 365 507
rect 541 779 542 781
rect 544 779 545 781
rect 541 785 542 787
rect 544 785 545 787
rect 561 119 562 121
rect 564 119 565 121
rect 561 125 562 127
rect 564 125 565 127
rect 741 619 742 621
rect 744 619 745 621
rect 741 625 742 627
rect 744 625 745 627
rect 541 359 542 361
rect 544 359 545 361
rect 541 365 542 367
rect 544 365 545 367
rect 321 439 322 441
rect 324 439 325 441
rect 321 445 322 447
rect 324 445 325 447
rect 661 459 662 461
rect 664 459 665 461
rect 661 465 662 467
rect 664 465 665 467
rect 581 239 582 241
rect 584 239 585 241
rect 581 245 582 247
rect 584 245 585 247
rect 461 819 462 821
rect 464 819 465 821
rect 461 825 462 827
rect 464 825 465 827
rect 621 739 622 741
rect 624 739 625 741
rect 621 745 622 747
rect 624 745 625 747
rect 661 659 662 661
rect 664 659 665 661
rect 661 665 662 667
rect 664 665 665 667
rect 501 319 502 321
rect 504 319 505 321
rect 501 325 502 327
rect 504 325 505 327
rect 701 459 702 461
rect 704 459 705 461
rect 701 465 702 467
rect 704 465 705 467
rect 661 599 662 601
rect 664 599 665 601
rect 661 605 662 607
rect 664 605 665 607
rect 441 699 442 701
rect 444 699 445 701
rect 441 705 442 707
rect 444 705 445 707
rect 241 319 242 321
rect 244 319 245 321
rect 241 325 242 327
rect 244 325 245 327
rect 321 659 322 661
rect 324 659 325 661
rect 321 665 322 667
rect 324 665 325 667
rect 361 719 362 721
rect 364 719 365 721
rect 361 725 362 727
rect 364 725 365 727
rect 401 659 402 661
rect 404 659 405 661
rect 401 665 402 667
rect 404 665 405 667
rect 641 819 642 821
rect 644 819 645 821
rect 641 825 642 827
rect 644 825 645 827
rect 241 699 242 701
rect 244 699 245 701
rect 241 705 242 707
rect 244 705 245 707
rect 621 799 622 801
rect 624 799 625 801
rect 621 805 622 807
rect 624 805 625 807
rect 261 479 262 481
rect 264 479 265 481
rect 261 485 262 487
rect 264 485 265 487
rect 741 459 742 461
rect 744 459 745 461
rect 741 465 742 467
rect 744 465 745 467
rect 681 699 682 701
rect 684 699 685 701
rect 681 705 682 707
rect 684 705 685 707
rect 521 719 522 721
rect 524 719 525 721
rect 521 725 522 727
rect 524 725 525 727
rect 601 339 602 341
rect 604 339 605 341
rect 601 345 602 347
rect 604 345 605 347
rect 441 859 442 861
rect 444 859 445 861
rect 441 865 442 867
rect 444 865 445 867
rect 561 479 562 481
rect 564 479 565 481
rect 561 485 562 487
rect 564 485 565 487
rect 681 259 682 261
rect 684 259 685 261
rect 681 265 682 267
rect 684 265 685 267
rect 481 399 482 401
rect 484 399 485 401
rect 481 405 482 407
rect 484 405 485 407
rect 721 459 722 461
rect 724 459 725 461
rect 721 465 722 467
rect 724 465 725 467
rect 381 239 382 241
rect 384 239 385 241
rect 381 245 382 247
rect 384 245 385 247
rect 441 679 442 681
rect 444 679 445 681
rect 441 685 442 687
rect 444 685 445 687
rect 401 739 402 741
rect 404 739 405 741
rect 401 745 402 747
rect 404 745 405 747
rect 641 419 642 421
rect 644 419 645 421
rect 641 425 642 427
rect 644 425 645 427
rect 281 519 282 521
rect 284 519 285 521
rect 281 525 282 527
rect 284 525 285 527
rect 701 559 702 561
rect 704 559 705 561
rect 701 565 702 567
rect 704 565 705 567
rect 341 619 342 621
rect 344 619 345 621
rect 341 625 342 627
rect 344 625 345 627
rect 521 439 522 441
rect 524 439 525 441
rect 521 445 522 447
rect 524 445 525 447
rect 541 159 542 161
rect 544 159 545 161
rect 541 165 542 167
rect 544 165 545 167
rect 441 339 442 341
rect 444 339 445 341
rect 441 345 442 347
rect 444 345 445 347
rect 801 559 802 561
rect 804 559 805 561
rect 801 565 802 567
rect 804 565 805 567
rect 481 819 482 821
rect 484 819 485 821
rect 481 825 482 827
rect 484 825 485 827
rect 241 619 242 621
rect 244 619 245 621
rect 241 625 242 627
rect 244 625 245 627
rect 321 779 322 781
rect 324 779 325 781
rect 321 785 322 787
rect 324 785 325 787
rect 361 619 362 621
rect 364 619 365 621
rect 361 625 362 627
rect 364 625 365 627
rect 701 759 702 761
rect 704 759 705 761
rect 701 765 702 767
rect 704 765 705 767
rect 421 579 422 581
rect 424 579 425 581
rect 421 585 422 587
rect 424 585 425 587
rect 681 659 682 661
rect 684 659 685 661
rect 681 665 682 667
rect 684 665 685 667
rect 321 259 322 261
rect 324 259 325 261
rect 321 265 322 267
rect 324 265 325 267
rect 801 419 802 421
rect 804 419 805 421
rect 801 425 802 427
rect 804 425 805 427
rect 321 459 322 461
rect 324 459 325 461
rect 321 465 322 467
rect 324 465 325 467
rect 701 359 702 361
rect 704 359 705 361
rect 701 365 702 367
rect 704 365 705 367
rect 601 559 602 561
rect 604 559 605 561
rect 601 565 602 567
rect 604 565 605 567
rect 241 579 242 581
rect 244 579 245 581
rect 241 585 242 587
rect 244 585 245 587
rect 741 639 742 641
rect 744 639 745 641
rect 741 645 742 647
rect 744 645 745 647
rect 741 399 742 401
rect 744 399 745 401
rect 741 405 742 407
rect 744 405 745 407
rect 661 219 662 221
rect 664 219 665 221
rect 661 225 662 227
rect 664 225 665 227
rect 101 519 102 521
rect 104 519 105 521
rect 101 525 102 527
rect 104 525 105 527
rect 361 519 362 521
rect 364 519 365 521
rect 361 525 362 527
rect 364 525 365 527
rect 421 319 422 321
rect 424 319 425 321
rect 421 325 422 327
rect 424 325 425 327
rect 501 719 502 721
rect 504 719 505 721
rect 501 725 502 727
rect 504 725 505 727
rect 741 379 742 381
rect 744 379 745 381
rect 741 385 742 387
rect 744 385 745 387
rect 221 679 222 681
rect 224 679 225 681
rect 221 685 222 687
rect 224 685 225 687
rect 421 359 422 361
rect 424 359 425 361
rect 421 365 422 367
rect 424 365 425 367
rect 261 519 262 521
rect 264 519 265 521
rect 261 525 262 527
rect 264 525 265 527
rect 781 419 782 421
rect 784 419 785 421
rect 781 425 782 427
rect 784 425 785 427
rect 381 639 382 641
rect 384 639 385 641
rect 381 645 382 647
rect 384 645 385 647
rect 521 539 522 541
rect 524 539 525 541
rect 521 545 522 547
rect 524 545 525 547
rect 721 579 722 581
rect 724 579 725 581
rect 721 585 722 587
rect 724 585 725 587
rect 441 459 442 461
rect 444 459 445 461
rect 441 465 442 467
rect 444 465 445 467
rect 661 379 662 381
rect 664 379 665 381
rect 661 385 662 387
rect 664 385 665 387
rect 421 259 422 261
rect 424 259 425 261
rect 421 265 422 267
rect 424 265 425 267
rect 521 699 522 701
rect 524 699 525 701
rect 521 705 522 707
rect 524 705 525 707
rect 681 479 682 481
rect 684 479 685 481
rect 681 485 682 487
rect 684 485 685 487
rect 681 439 682 441
rect 684 439 685 441
rect 681 445 682 447
rect 684 445 685 447
rect 361 559 362 561
rect 364 559 365 561
rect 361 565 362 567
rect 364 565 365 567
rect 601 219 602 221
rect 604 219 605 221
rect 601 225 602 227
rect 604 225 605 227
rect 521 779 522 781
rect 524 779 525 781
rect 521 785 522 787
rect 524 785 525 787
rect 261 679 262 681
rect 264 679 265 681
rect 261 685 262 687
rect 264 685 265 687
rect 541 439 542 441
rect 544 439 545 441
rect 541 445 542 447
rect 544 445 545 447
rect 321 699 322 701
rect 324 699 325 701
rect 321 705 322 707
rect 324 705 325 707
rect 761 379 762 381
rect 764 379 765 381
rect 761 385 762 387
rect 764 385 765 387
rect 421 659 422 661
rect 424 659 425 661
rect 421 665 422 667
rect 424 665 425 667
rect 221 439 222 441
rect 224 439 225 441
rect 221 445 222 447
rect 224 445 225 447
rect 361 419 362 421
rect 364 419 365 421
rect 361 425 362 427
rect 364 425 365 427
rect 781 659 782 661
rect 784 659 785 661
rect 781 665 782 667
rect 784 665 785 667
rect 461 799 462 801
rect 464 799 465 801
rect 461 805 462 807
rect 464 805 465 807
rect 721 659 722 661
rect 724 659 725 661
rect 721 665 722 667
rect 724 665 725 667
rect 561 359 562 361
rect 564 359 565 361
rect 561 365 562 367
rect 564 365 565 367
rect 601 279 602 281
rect 604 279 605 281
rect 601 285 602 287
rect 604 285 605 287
rect 381 459 382 461
rect 384 459 385 461
rect 381 465 382 467
rect 384 465 385 467
rect 581 399 582 401
rect 584 399 585 401
rect 581 405 582 407
rect 584 405 585 407
rect 521 259 522 261
rect 524 259 525 261
rect 521 265 522 267
rect 524 265 525 267
rect 621 299 622 301
rect 624 299 625 301
rect 621 305 622 307
rect 624 305 625 307
rect 281 459 282 461
rect 284 459 285 461
rect 281 465 282 467
rect 284 465 285 467
rect 301 439 302 441
rect 304 439 305 441
rect 301 445 302 447
rect 304 445 305 447
rect 501 199 502 201
rect 504 199 505 201
rect 501 205 502 207
rect 504 205 505 207
rect 141 639 142 641
rect 144 639 145 641
rect 141 645 142 647
rect 144 645 145 647
rect 641 619 642 621
rect 644 619 645 621
rect 641 625 642 627
rect 644 625 645 627
rect 401 339 402 341
rect 404 339 405 341
rect 401 345 402 347
rect 404 345 405 347
rect 881 539 882 541
rect 884 539 885 541
rect 881 545 882 547
rect 884 545 885 547
rect 761 519 762 521
rect 764 519 765 521
rect 761 525 762 527
rect 764 525 765 527
rect 421 459 422 461
rect 424 459 425 461
rect 421 465 422 467
rect 424 465 425 467
rect 481 419 482 421
rect 484 419 485 421
rect 481 425 482 427
rect 484 425 485 427
rect 521 839 522 841
rect 524 839 525 841
rect 521 845 522 847
rect 524 845 525 847
rect 541 659 542 661
rect 544 659 545 661
rect 541 665 542 667
rect 544 665 545 667
rect 461 599 462 601
rect 464 599 465 601
rect 461 605 462 607
rect 464 605 465 607
rect 461 499 462 501
rect 464 499 465 501
rect 461 505 462 507
rect 464 505 465 507
rect 781 499 782 501
rect 784 499 785 501
rect 781 505 782 507
rect 784 505 785 507
rect 341 759 342 761
rect 344 759 345 761
rect 341 765 342 767
rect 344 765 345 767
rect 261 399 262 401
rect 264 399 265 401
rect 261 405 262 407
rect 264 405 265 407
rect 441 279 442 281
rect 444 279 445 281
rect 441 285 442 287
rect 444 285 445 287
rect 681 179 682 181
rect 684 179 685 181
rect 681 185 682 187
rect 684 185 685 187
rect 221 499 222 501
rect 224 499 225 501
rect 221 505 222 507
rect 224 505 225 507
rect 621 839 622 841
rect 624 839 625 841
rect 621 845 622 847
rect 624 845 625 847
rect 541 239 542 241
rect 544 239 545 241
rect 541 245 542 247
rect 544 245 545 247
rect 361 379 362 381
rect 364 379 365 381
rect 361 385 362 387
rect 364 385 365 387
rect 721 479 722 481
rect 724 479 725 481
rect 721 485 722 487
rect 724 485 725 487
rect 281 619 282 621
rect 284 619 285 621
rect 281 625 282 627
rect 284 625 285 627
rect 241 339 242 341
rect 244 339 245 341
rect 241 345 242 347
rect 244 345 245 347
rect 361 739 362 741
rect 364 739 365 741
rect 361 745 362 747
rect 364 745 365 747
rect 381 319 382 321
rect 384 319 385 321
rect 381 325 382 327
rect 384 325 385 327
rect 381 379 382 381
rect 384 379 385 381
rect 381 385 382 387
rect 384 385 385 387
rect 201 579 202 581
rect 204 579 205 581
rect 201 585 202 587
rect 204 585 205 587
rect 401 239 402 241
rect 404 239 405 241
rect 401 245 402 247
rect 404 245 405 247
rect 241 559 242 561
rect 244 559 245 561
rect 241 565 242 567
rect 244 565 245 567
rect 721 519 722 521
rect 724 519 725 521
rect 721 525 722 527
rect 724 525 725 527
rect 661 639 662 641
rect 664 639 665 641
rect 661 645 662 647
rect 664 645 665 647
rect 301 599 302 601
rect 304 599 305 601
rect 301 605 302 607
rect 304 605 305 607
rect 501 739 502 741
rect 504 739 505 741
rect 501 745 502 747
rect 504 745 505 747
rect 601 199 602 201
rect 604 199 605 201
rect 601 205 602 207
rect 604 205 605 207
rect 581 879 582 881
rect 584 879 585 881
rect 581 885 582 887
rect 584 885 585 887
rect 181 499 182 501
rect 184 499 185 501
rect 181 505 182 507
rect 184 505 185 507
rect 581 659 582 661
rect 584 659 585 661
rect 581 665 582 667
rect 584 665 585 667
rect 661 439 662 441
rect 664 439 665 441
rect 661 445 662 447
rect 664 445 665 447
rect 521 459 522 461
rect 524 459 525 461
rect 521 465 522 467
rect 524 465 525 467
rect 461 739 462 741
rect 464 739 465 741
rect 461 745 462 747
rect 464 745 465 747
rect 441 199 442 201
rect 444 199 445 201
rect 441 205 442 207
rect 444 205 445 207
rect 861 559 862 561
rect 864 559 865 561
rect 861 565 862 567
rect 864 565 865 567
rect 301 299 302 301
rect 304 299 305 301
rect 301 305 302 307
rect 304 305 305 307
rect 301 659 302 661
rect 304 659 305 661
rect 301 665 302 667
rect 304 665 305 667
rect 761 399 762 401
rect 764 399 765 401
rect 761 405 762 407
rect 764 405 765 407
rect 341 479 342 481
rect 344 479 345 481
rect 341 485 342 487
rect 344 485 345 487
rect 481 179 482 181
rect 484 179 485 181
rect 481 185 482 187
rect 484 185 485 187
rect 241 519 242 521
rect 244 519 245 521
rect 241 525 242 527
rect 244 525 245 527
rect 641 719 642 721
rect 644 719 645 721
rect 641 725 642 727
rect 644 725 645 727
rect 441 319 442 321
rect 444 319 445 321
rect 441 325 442 327
rect 444 325 445 327
rect 801 539 802 541
rect 804 539 805 541
rect 801 545 802 547
rect 804 545 805 547
rect 341 539 342 541
rect 344 539 345 541
rect 341 545 342 547
rect 344 545 345 547
rect 541 279 542 281
rect 544 279 545 281
rect 541 285 542 287
rect 544 285 545 287
rect 701 399 702 401
rect 704 399 705 401
rect 701 405 702 407
rect 704 405 705 407
rect 541 579 542 581
rect 544 579 545 581
rect 541 585 542 587
rect 544 585 545 587
rect 321 799 322 801
rect 324 799 325 801
rect 321 805 322 807
rect 324 805 325 807
rect 341 499 342 501
rect 344 499 345 501
rect 341 505 342 507
rect 344 505 345 507
rect 541 679 542 681
rect 544 679 545 681
rect 541 685 542 687
rect 544 685 545 687
rect 561 699 562 701
rect 564 699 565 701
rect 561 705 562 707
rect 564 705 565 707
rect 721 299 722 301
rect 724 299 725 301
rect 721 305 722 307
rect 724 305 725 307
rect 561 219 562 221
rect 564 219 565 221
rect 561 225 562 227
rect 564 225 565 227
rect 421 219 422 221
rect 424 219 425 221
rect 421 225 422 227
rect 424 225 425 227
rect 521 219 522 221
rect 524 219 525 221
rect 521 225 522 227
rect 524 225 525 227
rect 281 379 282 381
rect 284 379 285 381
rect 281 385 282 387
rect 284 385 285 387
rect 761 419 762 421
rect 764 419 765 421
rect 761 425 762 427
rect 764 425 765 427
rect 501 539 502 541
rect 504 539 505 541
rect 501 545 502 547
rect 504 545 505 547
rect 441 559 442 561
rect 444 559 445 561
rect 441 565 442 567
rect 444 565 445 567
rect 521 619 522 621
rect 524 619 525 621
rect 521 625 522 627
rect 524 625 525 627
rect 121 519 122 521
rect 124 519 125 521
rect 121 525 122 527
rect 124 525 125 527
rect 601 699 602 701
rect 604 699 605 701
rect 601 705 602 707
rect 604 705 605 707
rect 881 479 882 481
rect 884 479 885 481
rect 881 485 882 487
rect 884 485 885 487
rect 641 459 642 461
rect 644 459 645 461
rect 641 465 642 467
rect 644 465 645 467
rect 501 819 502 821
rect 504 819 505 821
rect 501 825 502 827
rect 504 825 505 827
rect 501 459 502 461
rect 504 459 505 461
rect 501 465 502 467
rect 504 465 505 467
rect 301 579 302 581
rect 304 579 305 581
rect 301 585 302 587
rect 304 585 305 587
rect 641 279 642 281
rect 644 279 645 281
rect 641 285 642 287
rect 644 285 645 287
rect 401 319 402 321
rect 404 319 405 321
rect 401 325 402 327
rect 404 325 405 327
rect 281 319 282 321
rect 284 319 285 321
rect 281 325 282 327
rect 284 325 285 327
rect 801 359 802 361
rect 804 359 805 361
rect 801 365 802 367
rect 804 365 805 367
rect 621 679 622 681
rect 624 679 625 681
rect 621 685 622 687
rect 624 685 625 687
rect 521 199 522 201
rect 524 199 525 201
rect 521 205 522 207
rect 524 205 525 207
rect 841 559 842 561
rect 844 559 845 561
rect 841 565 842 567
rect 844 565 845 567
rect 441 579 442 581
rect 444 579 445 581
rect 441 585 442 587
rect 444 585 445 587
rect 501 619 502 621
rect 504 619 505 621
rect 501 625 502 627
rect 504 625 505 627
rect 501 559 502 561
rect 504 559 505 561
rect 501 565 502 567
rect 504 565 505 567
rect 281 559 282 561
rect 284 559 285 561
rect 281 565 282 567
rect 284 565 285 567
rect 481 739 482 741
rect 484 739 485 741
rect 481 745 482 747
rect 484 745 485 747
rect 641 399 642 401
rect 644 399 645 401
rect 641 405 642 407
rect 644 405 645 407
rect 581 259 582 261
rect 584 259 585 261
rect 581 265 582 267
rect 584 265 585 267
rect 221 519 222 521
rect 224 519 225 521
rect 221 525 222 527
rect 224 525 225 527
rect 401 779 402 781
rect 404 779 405 781
rect 401 785 402 787
rect 404 785 405 787
rect 501 239 502 241
rect 504 239 505 241
rect 501 245 502 247
rect 504 245 505 247
rect 721 559 722 561
rect 724 559 725 561
rect 721 565 722 567
rect 724 565 725 567
rect 421 179 422 181
rect 424 179 425 181
rect 421 185 422 187
rect 424 185 425 187
rect 241 499 242 501
rect 244 499 245 501
rect 241 505 242 507
rect 244 505 245 507
rect 581 439 582 441
rect 584 439 585 441
rect 581 445 582 447
rect 584 445 585 447
rect 781 519 782 521
rect 784 519 785 521
rect 781 525 782 527
rect 784 525 785 527
rect 681 679 682 681
rect 684 679 685 681
rect 681 685 682 687
rect 684 685 685 687
rect 261 639 262 641
rect 264 639 265 641
rect 261 645 262 647
rect 264 645 265 647
rect 861 519 862 521
rect 864 519 865 521
rect 861 525 862 527
rect 864 525 865 527
rect 541 419 542 421
rect 544 419 545 421
rect 541 425 542 427
rect 544 425 545 427
rect 521 159 522 161
rect 524 159 525 161
rect 521 165 522 167
rect 524 165 525 167
rect 561 879 562 881
rect 564 879 565 881
rect 561 885 562 887
rect 564 885 565 887
rect 321 419 322 421
rect 324 419 325 421
rect 321 425 322 427
rect 324 425 325 427
rect 541 519 542 521
rect 544 519 545 521
rect 541 525 542 527
rect 544 525 545 527
rect 581 719 582 721
rect 584 719 585 721
rect 581 725 582 727
rect 584 725 585 727
rect 201 679 202 681
rect 204 679 205 681
rect 201 685 202 687
rect 204 685 205 687
rect 361 579 362 581
rect 364 579 365 581
rect 361 585 362 587
rect 364 585 365 587
rect 621 399 622 401
rect 624 399 625 401
rect 621 405 622 407
rect 624 405 625 407
rect 561 399 562 401
rect 564 399 565 401
rect 561 405 562 407
rect 564 405 565 407
rect 561 259 562 261
rect 564 259 565 261
rect 561 265 562 267
rect 564 265 565 267
rect 761 599 762 601
rect 764 599 765 601
rect 761 605 762 607
rect 764 605 765 607
rect 481 259 482 261
rect 484 259 485 261
rect 481 265 482 267
rect 484 265 485 267
rect 621 759 622 761
rect 624 759 625 761
rect 621 765 622 767
rect 624 765 625 767
rect 761 459 762 461
rect 764 459 765 461
rect 761 465 762 467
rect 764 465 765 467
rect 621 559 622 561
rect 624 559 625 561
rect 621 565 622 567
rect 624 565 625 567
rect 781 699 782 701
rect 784 699 785 701
rect 781 705 782 707
rect 784 705 785 707
rect 581 579 582 581
rect 584 579 585 581
rect 581 585 582 587
rect 584 585 585 587
rect 461 579 462 581
rect 464 579 465 581
rect 461 585 462 587
rect 464 585 465 587
rect 581 419 582 421
rect 584 419 585 421
rect 581 425 582 427
rect 584 425 585 427
rect 661 779 662 781
rect 664 779 665 781
rect 661 785 662 787
rect 664 785 665 787
rect 821 439 822 441
rect 824 439 825 441
rect 821 445 822 447
rect 824 445 825 447
rect 501 279 502 281
rect 504 279 505 281
rect 501 285 502 287
rect 504 285 505 287
rect 561 459 562 461
rect 564 459 565 461
rect 561 465 562 467
rect 564 465 565 467
rect 161 399 162 401
rect 164 399 165 401
rect 161 405 162 407
rect 164 405 165 407
rect 581 559 582 561
rect 584 559 585 561
rect 581 565 582 567
rect 584 565 585 567
rect 581 699 582 701
rect 584 699 585 701
rect 581 705 582 707
rect 584 705 585 707
rect 821 499 822 501
rect 824 499 825 501
rect 821 505 822 507
rect 824 505 825 507
rect 721 739 722 741
rect 724 739 725 741
rect 721 745 722 747
rect 724 745 725 747
rect 441 759 442 761
rect 444 759 445 761
rect 441 765 442 767
rect 444 765 445 767
rect 761 319 762 321
rect 764 319 765 321
rect 761 325 762 327
rect 764 325 765 327
rect 341 699 342 701
rect 344 699 345 701
rect 341 705 342 707
rect 344 705 345 707
rect 721 359 722 361
rect 724 359 725 361
rect 721 365 722 367
rect 724 365 725 367
rect 701 699 702 701
rect 704 699 705 701
rect 701 705 702 707
rect 704 705 705 707
rect 521 759 522 761
rect 524 759 525 761
rect 521 765 522 767
rect 524 765 525 767
rect 521 359 522 361
rect 524 359 525 361
rect 521 365 522 367
rect 524 365 525 367
rect 421 559 422 561
rect 424 559 425 561
rect 421 565 422 567
rect 424 565 425 567
rect 161 539 162 541
rect 164 539 165 541
rect 161 545 162 547
rect 164 545 165 547
rect 341 679 342 681
rect 344 679 345 681
rect 341 685 342 687
rect 344 685 345 687
rect 681 359 682 361
rect 684 359 685 361
rect 681 365 682 367
rect 684 365 685 367
rect 221 659 222 661
rect 224 659 225 661
rect 221 665 222 667
rect 224 665 225 667
rect 141 499 142 501
rect 144 499 145 501
rect 141 505 142 507
rect 144 505 145 507
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
rect -19 -21 -18 -19
rect -16 -21 -15 -19
rect -19 -15 -18 -13
rect -16 -15 -15 -13
<< labels >>
rlabel pdiffusion 363 263 364 264 0 Cellno = 1
rlabel pdiffusion 723 423 724 424 0 Cellno = 2
rlabel pdiffusion 203 383 204 384 0 Cellno = 3
rlabel pdiffusion 743 483 744 484 0 Cellno = 4
rlabel pdiffusion 623 823 624 824 0 Cellno = 5
rlabel pdiffusion 263 543 264 544 0 Cellno = 6
rlabel pdiffusion 383 403 384 404 0 Cellno = 7
rlabel pdiffusion 503 423 504 424 0 Cellno = 8
rlabel pdiffusion 263 363 264 364 0 Cellno = 9
rlabel pdiffusion 263 663 264 664 0 Cellno = 10
rlabel pdiffusion 763 663 764 664 0 Cellno = 11
rlabel pdiffusion 383 663 384 664 0 Cellno = 12
rlabel pdiffusion 483 803 484 804 0 Cellno = 13
rlabel pdiffusion 743 683 744 684 0 Cellno = 14
rlabel pdiffusion 183 483 184 484 0 Cellno = 15
rlabel pdiffusion 603 623 604 624 0 Cellno = 16
rlabel pdiffusion 863 543 864 544 0 Cellno = 17
rlabel pdiffusion 563 583 564 584 0 Cellno = 18
rlabel pdiffusion 663 623 664 624 0 Cellno = 19
rlabel pdiffusion 323 383 324 384 0 Cellno = 20
rlabel pdiffusion 583 803 584 804 0 Cellno = 21
rlabel pdiffusion 203 443 204 444 0 Cellno = 22
rlabel pdiffusion 323 583 324 584 0 Cellno = 23
rlabel pdiffusion 223 363 224 364 0 Cellno = 24
rlabel pdiffusion 263 343 264 344 0 Cellno = 25
rlabel pdiffusion 643 563 644 564 0 Cellno = 26
rlabel pdiffusion 163 443 164 444 0 Cellno = 27
rlabel pdiffusion 623 723 624 724 0 Cellno = 28
rlabel pdiffusion 463 723 464 724 0 Cellno = 29
rlabel pdiffusion 483 663 484 664 0 Cellno = 30
rlabel pdiffusion 603 463 604 464 0 Cellno = 31
rlabel pdiffusion 383 483 384 484 0 Cellno = 32
rlabel pdiffusion 723 683 724 684 0 Cellno = 33
rlabel pdiffusion 543 463 544 464 0 Cellno = 34
rlabel pdiffusion 623 503 624 504 0 Cellno = 35
rlabel pdiffusion 383 283 384 284 0 Cellno = 36
rlabel pdiffusion 823 663 824 664 0 Cellno = 37
rlabel pdiffusion 123 503 124 504 0 Cellno = 38
rlabel pdiffusion 503 803 504 804 0 Cellno = 39
rlabel pdiffusion 643 303 644 304 0 Cellno = 40
rlabel pdiffusion 803 463 804 464 0 Cellno = 41
rlabel pdiffusion 483 283 484 284 0 Cellno = 42
rlabel pdiffusion 743 703 744 704 0 Cellno = 43
rlabel pdiffusion 803 383 804 384 0 Cellno = 44
rlabel pdiffusion 423 683 424 684 0 Cellno = 45
rlabel pdiffusion 443 183 444 184 0 Cellno = 46
rlabel pdiffusion 503 843 504 844 0 Cellno = 47
rlabel pdiffusion 543 643 544 644 0 Cellno = 48
rlabel pdiffusion 623 263 624 264 0 Cellno = 49
rlabel pdiffusion 483 863 484 864 0 Cellno = 50
rlabel pdiffusion 443 803 444 804 0 Cellno = 51
rlabel pdiffusion 823 463 824 464 0 Cellno = 52
rlabel pdiffusion 603 743 604 744 0 Cellno = 53
rlabel pdiffusion 463 683 464 684 0 Cellno = 54
rlabel pdiffusion 223 483 224 484 0 Cellno = 55
rlabel pdiffusion 663 543 664 544 0 Cellno = 56
rlabel pdiffusion 343 723 344 724 0 Cellno = 57
rlabel pdiffusion 443 883 444 884 0 Cellno = 58
rlabel pdiffusion 403 803 404 804 0 Cellno = 59
rlabel pdiffusion 143 583 144 584 0 Cellno = 60
rlabel pdiffusion 183 583 184 584 0 Cellno = 61
rlabel pdiffusion 723 723 724 724 0 Cellno = 62
rlabel pdiffusion 323 483 324 484 0 Cellno = 63
rlabel pdiffusion 623 623 624 624 0 Cellno = 64
rlabel pdiffusion 563 803 564 804 0 Cellno = 65
rlabel pdiffusion 283 763 284 764 0 Cellno = 66
rlabel pdiffusion 803 683 804 684 0 Cellno = 67
rlabel pdiffusion 543 563 544 564 0 Cellno = 68
rlabel pdiffusion 443 503 444 504 0 Cellno = 69
rlabel pdiffusion 783 383 784 384 0 Cellno = 70
rlabel pdiffusion 803 603 804 604 0 Cellno = 71
rlabel pdiffusion 643 703 644 704 0 Cellno = 72
rlabel pdiffusion 503 763 504 764 0 Cellno = 73
rlabel pdiffusion 323 363 324 364 0 Cellno = 74
rlabel pdiffusion 163 563 164 564 0 Cellno = 75
rlabel pdiffusion 423 383 424 384 0 Cellno = 76
rlabel pdiffusion 143 623 144 624 0 Cellno = 77
rlabel pdiffusion 683 583 684 584 0 Cellno = 78
rlabel pdiffusion 783 623 784 624 0 Cellno = 79
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 80
rlabel pdiffusion 323 623 324 624 0 Cellno = 81
rlabel pdiffusion 723 443 724 444 0 Cellno = 82
rlabel pdiffusion 483 583 484 584 0 Cellno = 83
rlabel pdiffusion 343 743 344 744 0 Cellno = 84
rlabel pdiffusion 183 643 184 644 0 Cellno = 85
rlabel pdiffusion 803 443 804 444 0 Cellno = 86
rlabel pdiffusion 663 323 664 324 0 Cellno = 87
rlabel pdiffusion 263 743 264 744 0 Cellno = 88
rlabel pdiffusion 383 203 384 204 0 Cellno = 89
rlabel pdiffusion 623 383 624 384 0 Cellno = 90
rlabel pdiffusion 643 803 644 804 0 Cellno = 91
rlabel pdiffusion 483 163 484 164 0 Cellno = 92
rlabel pdiffusion 263 723 264 724 0 Cellno = 93
rlabel pdiffusion 583 483 584 484 0 Cellno = 94
rlabel pdiffusion 443 783 444 784 0 Cellno = 95
rlabel pdiffusion 863 503 864 504 0 Cellno = 96
rlabel pdiffusion 843 403 844 404 0 Cellno = 97
rlabel pdiffusion 323 603 324 604 0 Cellno = 98
rlabel pdiffusion 523 823 524 824 0 Cellno = 99
rlabel pdiffusion 523 863 524 864 0 Cellno = 100
rlabel pdiffusion 483 643 484 644 0 Cellno = 101
rlabel pdiffusion 723 503 724 504 0 Cellno = 102
rlabel pdiffusion 663 203 664 204 0 Cellno = 103
rlabel pdiffusion 403 423 404 424 0 Cellno = 104
rlabel pdiffusion 403 823 404 824 0 Cellno = 105
rlabel pdiffusion 743 303 744 304 0 Cellno = 106
rlabel pdiffusion 463 623 464 624 0 Cellno = 107
rlabel pdiffusion 623 703 624 704 0 Cellno = 108
rlabel pdiffusion 163 583 164 584 0 Cellno = 109
rlabel pdiffusion 463 663 464 664 0 Cellno = 110
rlabel pdiffusion 263 383 264 384 0 Cellno = 111
rlabel pdiffusion 563 643 564 644 0 Cellno = 112
rlabel pdiffusion 343 443 344 444 0 Cellno = 113
rlabel pdiffusion 283 303 284 304 0 Cellno = 114
rlabel pdiffusion 403 263 404 264 0 Cellno = 115
rlabel pdiffusion 503 863 504 864 0 Cellno = 116
rlabel pdiffusion 403 223 404 224 0 Cellno = 117
rlabel pdiffusion 363 223 364 224 0 Cellno = 118
rlabel pdiffusion 763 483 764 484 0 Cellno = 119
rlabel pdiffusion 643 503 644 504 0 Cellno = 120
rlabel pdiffusion 523 583 524 584 0 Cellno = 121
rlabel pdiffusion 383 523 384 524 0 Cellno = 122
rlabel pdiffusion 463 443 464 444 0 Cellno = 123
rlabel pdiffusion 783 363 784 364 0 Cellno = 124
rlabel pdiffusion 543 903 544 904 0 Cellno = 125
rlabel pdiffusion 363 803 364 804 0 Cellno = 126
rlabel pdiffusion 183 543 184 544 0 Cellno = 127
rlabel pdiffusion 263 503 264 504 0 Cellno = 128
rlabel pdiffusion 383 723 384 724 0 Cellno = 129
rlabel pdiffusion 483 303 484 304 0 Cellno = 130
rlabel pdiffusion 303 383 304 384 0 Cellno = 131
rlabel pdiffusion 423 203 424 204 0 Cellno = 132
rlabel pdiffusion 583 203 584 204 0 Cellno = 133
rlabel pdiffusion 563 663 564 664 0 Cellno = 134
rlabel pdiffusion 643 843 644 844 0 Cellno = 135
rlabel pdiffusion 423 603 424 604 0 Cellno = 136
rlabel pdiffusion 283 503 284 504 0 Cellno = 137
rlabel pdiffusion 423 403 424 404 0 Cellno = 138
rlabel pdiffusion 683 403 684 404 0 Cellno = 139
rlabel pdiffusion 243 383 244 384 0 Cellno = 140
rlabel pdiffusion 323 643 324 644 0 Cellno = 141
rlabel pdiffusion 323 343 324 344 0 Cellno = 142
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 143
rlabel pdiffusion 403 543 404 544 0 Cellno = 144
rlabel pdiffusion 303 483 304 484 0 Cellno = 145
rlabel pdiffusion 423 343 424 344 0 Cellno = 146
rlabel pdiffusion 823 523 824 524 0 Cellno = 147
rlabel pdiffusion 203 663 204 664 0 Cellno = 148
rlabel pdiffusion 603 423 604 424 0 Cellno = 149
rlabel pdiffusion 823 583 824 584 0 Cellno = 150
rlabel pdiffusion 363 343 364 344 0 Cellno = 151
rlabel pdiffusion 643 543 644 544 0 Cellno = 152
rlabel pdiffusion 643 343 644 344 0 Cellno = 153
rlabel pdiffusion 483 463 484 464 0 Cellno = 154
rlabel pdiffusion 483 343 484 344 0 Cellno = 155
rlabel pdiffusion 363 443 364 444 0 Cellno = 156
rlabel pdiffusion 663 343 664 344 0 Cellno = 157
rlabel pdiffusion 283 743 284 744 0 Cellno = 158
rlabel pdiffusion 703 503 704 504 0 Cellno = 159
rlabel pdiffusion 263 323 264 324 0 Cellno = 160
rlabel pdiffusion 383 343 384 344 0 Cellno = 161
rlabel pdiffusion 703 543 704 544 0 Cellno = 162
rlabel pdiffusion 883 523 884 524 0 Cellno = 163
rlabel pdiffusion 843 543 844 544 0 Cellno = 164
rlabel pdiffusion 623 783 624 784 0 Cellno = 165
rlabel pdiffusion 323 543 324 544 0 Cellno = 166
rlabel pdiffusion 763 703 764 704 0 Cellno = 167
rlabel pdiffusion 363 783 364 784 0 Cellno = 168
rlabel pdiffusion 423 823 424 824 0 Cellno = 169
rlabel pdiffusion 743 723 744 724 0 Cellno = 170
rlabel pdiffusion 683 603 684 604 0 Cellno = 171
rlabel pdiffusion 643 223 644 224 0 Cellno = 172
rlabel pdiffusion 643 323 644 324 0 Cellno = 173
rlabel pdiffusion 783 643 784 644 0 Cellno = 174
rlabel pdiffusion 803 623 804 624 0 Cellno = 175
rlabel pdiffusion 463 223 464 224 0 Cellno = 176
rlabel pdiffusion 503 523 504 524 0 Cellno = 177
rlabel pdiffusion 443 303 444 304 0 Cellno = 178
rlabel pdiffusion 103 463 104 464 0 Cellno = 179
rlabel pdiffusion 183 523 184 524 0 Cellno = 180
rlabel pdiffusion 263 563 264 564 0 Cellno = 181
rlabel pdiffusion 603 403 604 404 0 Cellno = 182
rlabel pdiffusion 523 663 524 664 0 Cellno = 183
rlabel pdiffusion 143 523 144 524 0 Cellno = 184
rlabel pdiffusion 803 403 804 404 0 Cellno = 185
rlabel pdiffusion 583 823 584 824 0 Cellno = 186
rlabel pdiffusion 563 543 564 544 0 Cellno = 187
rlabel pdiffusion 203 503 204 504 0 Cellno = 188
rlabel pdiffusion 703 343 704 344 0 Cellno = 189
rlabel pdiffusion 563 423 564 424 0 Cellno = 190
rlabel pdiffusion 143 603 144 604 0 Cellno = 191
rlabel pdiffusion 503 383 504 384 0 Cellno = 192
rlabel pdiffusion 603 803 604 804 0 Cellno = 193
rlabel pdiffusion 443 623 444 624 0 Cellno = 194
rlabel pdiffusion 203 543 204 544 0 Cellno = 195
rlabel pdiffusion 163 423 164 424 0 Cellno = 196
rlabel pdiffusion 563 163 564 164 0 Cellno = 197
rlabel pdiffusion 383 763 384 764 0 Cellno = 198
rlabel pdiffusion 903 563 904 564 0 Cellno = 199
rlabel pdiffusion 283 603 284 604 0 Cellno = 200
rlabel pdiffusion 523 523 524 524 0 Cellno = 201
rlabel pdiffusion 523 423 524 424 0 Cellno = 202
rlabel pdiffusion 343 263 344 264 0 Cellno = 203
rlabel pdiffusion 203 523 204 524 0 Cellno = 204
rlabel pdiffusion 763 503 764 504 0 Cellno = 205
rlabel pdiffusion 883 503 884 504 0 Cellno = 206
rlabel pdiffusion 363 763 364 764 0 Cellno = 207
rlabel pdiffusion 583 783 584 784 0 Cellno = 208
rlabel pdiffusion 623 183 624 184 0 Cellno = 209
rlabel pdiffusion 343 403 344 404 0 Cellno = 210
rlabel pdiffusion 443 543 444 544 0 Cellno = 211
rlabel pdiffusion 823 603 824 604 0 Cellno = 212
rlabel pdiffusion 363 283 364 284 0 Cellno = 213
rlabel pdiffusion 543 503 544 504 0 Cellno = 214
rlabel pdiffusion 543 183 544 184 0 Cellno = 215
rlabel pdiffusion 403 763 404 764 0 Cellno = 216
rlabel pdiffusion 703 303 704 304 0 Cellno = 217
rlabel pdiffusion 283 543 284 544 0 Cellno = 218
rlabel pdiffusion 783 683 784 684 0 Cellno = 219
rlabel pdiffusion 183 663 184 664 0 Cellno = 220
rlabel pdiffusion 443 243 444 244 0 Cellno = 221
rlabel pdiffusion 343 823 344 824 0 Cellno = 222
rlabel pdiffusion 583 323 584 324 0 Cellno = 223
rlabel pdiffusion 323 723 324 724 0 Cellno = 224
rlabel pdiffusion 503 583 504 584 0 Cellno = 225
rlabel pdiffusion 543 143 544 144 0 Cellno = 226
rlabel pdiffusion 403 563 404 564 0 Cellno = 227
rlabel pdiffusion 663 503 664 504 0 Cellno = 228
rlabel pdiffusion 203 623 204 624 0 Cellno = 229
rlabel pdiffusion 583 763 584 764 0 Cellno = 230
rlabel pdiffusion 123 443 124 444 0 Cellno = 231
rlabel pdiffusion 483 843 484 844 0 Cellno = 232
rlabel pdiffusion 483 763 484 764 0 Cellno = 233
rlabel pdiffusion 303 423 304 424 0 Cellno = 234
rlabel pdiffusion 823 643 824 644 0 Cellno = 235
rlabel pdiffusion 523 563 524 564 0 Cellno = 236
rlabel pdiffusion 503 883 504 884 0 Cellno = 237
rlabel pdiffusion 323 503 324 504 0 Cellno = 238
rlabel pdiffusion 883 463 884 464 0 Cellno = 239
rlabel pdiffusion 583 223 584 224 0 Cellno = 240
rlabel pdiffusion 803 643 804 644 0 Cellno = 241
rlabel pdiffusion 163 523 164 524 0 Cellno = 242
rlabel pdiffusion 643 583 644 584 0 Cellno = 243
rlabel pdiffusion 543 323 544 324 0 Cellno = 244
rlabel pdiffusion 283 443 284 444 0 Cellno = 245
rlabel pdiffusion 603 843 604 844 0 Cellno = 246
rlabel pdiffusion 803 503 804 504 0 Cellno = 247
rlabel pdiffusion 303 723 304 724 0 Cellno = 248
rlabel pdiffusion 683 523 684 524 0 Cellno = 249
rlabel pdiffusion 423 843 424 844 0 Cellno = 250
rlabel pdiffusion 403 443 404 444 0 Cellno = 251
rlabel pdiffusion 443 363 444 364 0 Cellno = 252
rlabel pdiffusion 843 463 844 464 0 Cellno = 253
rlabel pdiffusion 303 743 304 744 0 Cellno = 254
rlabel pdiffusion 283 723 284 724 0 Cellno = 255
rlabel pdiffusion 383 603 384 604 0 Cellno = 256
rlabel pdiffusion 603 823 604 824 0 Cellno = 257
rlabel pdiffusion 483 323 484 324 0 Cellno = 258
rlabel pdiffusion 743 443 744 444 0 Cellno = 259
rlabel pdiffusion 483 543 484 544 0 Cellno = 260
rlabel pdiffusion 543 843 544 844 0 Cellno = 261
rlabel pdiffusion 443 843 444 844 0 Cellno = 262
rlabel pdiffusion 463 863 464 864 0 Cellno = 263
rlabel pdiffusion 303 703 304 704 0 Cellno = 264
rlabel pdiffusion 463 523 464 524 0 Cellno = 265
rlabel pdiffusion 423 803 424 804 0 Cellno = 266
rlabel pdiffusion 523 603 524 604 0 Cellno = 267
rlabel pdiffusion 763 723 764 724 0 Cellno = 268
rlabel pdiffusion 343 563 344 564 0 Cellno = 269
rlabel pdiffusion 503 183 504 184 0 Cellno = 270
rlabel pdiffusion 443 383 444 384 0 Cellno = 271
rlabel pdiffusion 283 343 284 344 0 Cellno = 272
rlabel pdiffusion 223 563 224 564 0 Cellno = 273
rlabel pdiffusion 843 443 844 444 0 Cellno = 274
rlabel pdiffusion 243 683 244 684 0 Cellno = 275
rlabel pdiffusion 503 603 504 604 0 Cellno = 276
rlabel pdiffusion 743 743 744 744 0 Cellno = 277
rlabel pdiffusion 203 363 204 364 0 Cellno = 278
rlabel pdiffusion 163 623 164 624 0 Cellno = 279
rlabel pdiffusion 283 583 284 584 0 Cellno = 280
rlabel pdiffusion 743 603 744 604 0 Cellno = 281
rlabel pdiffusion 463 843 464 844 0 Cellno = 282
rlabel pdiffusion 683 383 684 384 0 Cellno = 283
rlabel pdiffusion 243 443 244 444 0 Cellno = 284
rlabel pdiffusion 643 783 644 784 0 Cellno = 285
rlabel pdiffusion 463 343 464 344 0 Cellno = 286
rlabel pdiffusion 743 663 744 664 0 Cellno = 287
rlabel pdiffusion 363 603 364 604 0 Cellno = 288
rlabel pdiffusion 423 483 424 484 0 Cellno = 289
rlabel pdiffusion 703 663 704 664 0 Cellno = 290
rlabel pdiffusion 343 323 344 324 0 Cellno = 291
rlabel pdiffusion 543 543 544 544 0 Cellno = 292
rlabel pdiffusion 223 463 224 464 0 Cellno = 293
rlabel pdiffusion 863 463 864 464 0 Cellno = 294
rlabel pdiffusion 563 743 564 744 0 Cellno = 295
rlabel pdiffusion 163 603 164 604 0 Cellno = 296
rlabel pdiffusion 643 263 644 264 0 Cellno = 297
rlabel pdiffusion 723 263 724 264 0 Cellno = 298
rlabel pdiffusion 783 543 784 544 0 Cellno = 299
rlabel pdiffusion 563 723 564 724 0 Cellno = 300
rlabel pdiffusion 503 263 504 264 0 Cellno = 301
rlabel pdiffusion 243 643 244 644 0 Cellno = 302
rlabel pdiffusion 463 403 464 404 0 Cellno = 303
rlabel pdiffusion 743 323 744 324 0 Cellno = 304
rlabel pdiffusion 363 703 364 704 0 Cellno = 305
rlabel pdiffusion 443 723 444 724 0 Cellno = 306
rlabel pdiffusion 403 623 404 624 0 Cellno = 307
rlabel pdiffusion 423 423 424 424 0 Cellno = 308
rlabel pdiffusion 223 403 224 404 0 Cellno = 309
rlabel pdiffusion 743 583 744 584 0 Cellno = 310
rlabel pdiffusion 463 263 464 264 0 Cellno = 311
rlabel pdiffusion 743 523 744 524 0 Cellno = 312
rlabel pdiffusion 463 783 464 784 0 Cellno = 313
rlabel pdiffusion 103 563 104 564 0 Cellno = 314
rlabel pdiffusion 483 723 484 724 0 Cellno = 315
rlabel pdiffusion 583 683 584 684 0 Cellno = 316
rlabel pdiffusion 543 763 544 764 0 Cellno = 317
rlabel pdiffusion 423 283 424 284 0 Cellno = 318
rlabel pdiffusion 683 243 684 244 0 Cellno = 319
rlabel pdiffusion 163 503 164 504 0 Cellno = 320
rlabel pdiffusion 643 523 644 524 0 Cellno = 321
rlabel pdiffusion 863 483 864 484 0 Cellno = 322
rlabel pdiffusion 683 723 684 724 0 Cellno = 323
rlabel pdiffusion 463 183 464 184 0 Cellno = 324
rlabel pdiffusion 563 863 564 864 0 Cellno = 325
rlabel pdiffusion 243 363 244 364 0 Cellno = 326
rlabel pdiffusion 703 283 704 284 0 Cellno = 327
rlabel pdiffusion 263 703 264 704 0 Cellno = 328
rlabel pdiffusion 143 443 144 444 0 Cellno = 329
rlabel pdiffusion 243 543 244 544 0 Cellno = 330
rlabel pdiffusion 843 623 844 624 0 Cellno = 331
rlabel pdiffusion 783 343 784 344 0 Cellno = 332
rlabel pdiffusion 223 423 224 424 0 Cellno = 333
rlabel pdiffusion 563 283 564 284 0 Cellno = 334
rlabel pdiffusion 463 423 464 424 0 Cellno = 335
rlabel pdiffusion 423 703 424 704 0 Cellno = 336
rlabel pdiffusion 143 563 144 564 0 Cellno = 337
rlabel pdiffusion 683 503 684 504 0 Cellno = 338
rlabel pdiffusion 823 563 824 564 0 Cellno = 339
rlabel pdiffusion 563 323 564 324 0 Cellno = 340
rlabel pdiffusion 843 583 844 584 0 Cellno = 341
rlabel pdiffusion 563 763 564 764 0 Cellno = 342
rlabel pdiffusion 703 683 704 684 0 Cellno = 343
rlabel pdiffusion 443 603 444 604 0 Cellno = 344
rlabel pdiffusion 503 783 504 784 0 Cellno = 345
rlabel pdiffusion 503 223 504 224 0 Cellno = 346
rlabel pdiffusion 263 463 264 464 0 Cellno = 347
rlabel pdiffusion 543 263 544 264 0 Cellno = 348
rlabel pdiffusion 663 283 664 284 0 Cellno = 349
rlabel pdiffusion 623 223 624 224 0 Cellno = 350
rlabel pdiffusion 723 283 724 284 0 Cellno = 351
rlabel pdiffusion 683 563 684 564 0 Cellno = 352
rlabel pdiffusion 703 623 704 624 0 Cellno = 353
rlabel pdiffusion 823 783 824 784 0 Cellno = 354
rlabel pdiffusion 243 423 244 424 0 Cellno = 355
rlabel pdiffusion 343 303 344 304 0 Cellno = 356
rlabel pdiffusion 583 163 584 164 0 Cellno = 357
rlabel pdiffusion 503 683 504 684 0 Cellno = 358
rlabel pdiffusion 823 403 824 404 0 Cellno = 359
rlabel pdiffusion 423 503 424 504 0 Cellno = 360
rlabel pdiffusion 703 423 704 424 0 Cellno = 361
rlabel pdiffusion 623 203 624 204 0 Cellno = 362
rlabel pdiffusion 483 223 484 224 0 Cellno = 363
rlabel pdiffusion 143 543 144 544 0 Cellno = 364
rlabel pdiffusion 243 663 244 664 0 Cellno = 365
rlabel pdiffusion 543 203 544 204 0 Cellno = 366
rlabel pdiffusion 383 423 384 424 0 Cellno = 367
rlabel pdiffusion 443 823 444 824 0 Cellno = 368
rlabel pdiffusion 283 403 284 404 0 Cellno = 369
rlabel pdiffusion 663 243 664 244 0 Cellno = 370
rlabel pdiffusion 223 603 224 604 0 Cellno = 371
rlabel pdiffusion 463 303 464 304 0 Cellno = 372
rlabel pdiffusion 183 423 184 424 0 Cellno = 373
rlabel pdiffusion 383 263 384 264 0 Cellno = 374
rlabel pdiffusion 303 323 304 324 0 Cellno = 375
rlabel pdiffusion 183 563 184 564 0 Cellno = 376
rlabel pdiffusion 383 683 384 684 0 Cellno = 377
rlabel pdiffusion 843 503 844 504 0 Cellno = 378
rlabel pdiffusion 463 643 464 644 0 Cellno = 379
rlabel pdiffusion 523 643 524 644 0 Cellno = 380
rlabel pdiffusion 763 363 764 364 0 Cellno = 381
rlabel pdiffusion 343 783 344 784 0 Cellno = 382
rlabel pdiffusion 623 443 624 444 0 Cellno = 383
rlabel pdiffusion 523 283 524 284 0 Cellno = 384
rlabel pdiffusion 503 403 504 404 0 Cellno = 385
rlabel pdiffusion 343 583 344 584 0 Cellno = 386
rlabel pdiffusion 823 483 824 484 0 Cellno = 387
rlabel pdiffusion 543 483 544 484 0 Cellno = 388
rlabel pdiffusion 343 383 344 384 0 Cellno = 389
rlabel pdiffusion 463 463 464 464 0 Cellno = 390
rlabel pdiffusion 563 243 564 244 0 Cellno = 391
rlabel pdiffusion 603 783 604 784 0 Cellno = 392
rlabel pdiffusion 503 663 504 664 0 Cellno = 393
rlabel pdiffusion 283 483 284 484 0 Cellno = 394
rlabel pdiffusion 783 443 784 444 0 Cellno = 395
rlabel pdiffusion 483 243 484 244 0 Cellno = 396
rlabel pdiffusion 703 743 704 744 0 Cellno = 397
rlabel pdiffusion 543 403 544 404 0 Cellno = 398
rlabel pdiffusion 443 163 444 164 0 Cellno = 399
rlabel pdiffusion 123 603 124 604 0 Cellno = 400
rlabel pdiffusion 703 583 704 584 0 Cellno = 401
rlabel pdiffusion 463 543 464 544 0 Cellno = 402
rlabel pdiffusion 403 303 404 304 0 Cellno = 403
rlabel pdiffusion 323 323 324 324 0 Cellno = 404
rlabel pdiffusion 263 583 264 584 0 Cellno = 405
rlabel pdiffusion 563 603 564 604 0 Cellno = 406
rlabel pdiffusion 643 183 644 184 0 Cellno = 407
rlabel pdiffusion 723 763 724 764 0 Cellno = 408
rlabel pdiffusion 123 463 124 464 0 Cellno = 409
rlabel pdiffusion 403 603 404 604 0 Cellno = 410
rlabel pdiffusion 523 403 524 404 0 Cellno = 411
rlabel pdiffusion 683 203 684 204 0 Cellno = 412
rlabel pdiffusion 623 523 624 524 0 Cellno = 413
rlabel pdiffusion 263 603 264 604 0 Cellno = 414
rlabel pdiffusion 523 743 524 744 0 Cellno = 415
rlabel pdiffusion 623 423 624 424 0 Cellno = 416
rlabel pdiffusion 283 683 284 684 0 Cellno = 417
rlabel pdiffusion 423 643 424 644 0 Cellno = 418
rlabel pdiffusion 563 303 564 304 0 Cellno = 419
rlabel pdiffusion 323 683 324 684 0 Cellno = 420
rlabel pdiffusion 563 503 564 504 0 Cellno = 421
rlabel pdiffusion 243 483 244 484 0 Cellno = 422
rlabel pdiffusion 703 603 704 604 0 Cellno = 423
rlabel pdiffusion 283 643 284 644 0 Cellno = 424
rlabel pdiffusion 303 563 304 564 0 Cellno = 425
rlabel pdiffusion 443 443 444 444 0 Cellno = 426
rlabel pdiffusion 603 443 604 444 0 Cellno = 427
rlabel pdiffusion 623 463 624 464 0 Cellno = 428
rlabel pdiffusion 663 583 664 584 0 Cellno = 429
rlabel pdiffusion 403 643 404 644 0 Cellno = 430
rlabel pdiffusion 263 443 264 444 0 Cellno = 431
rlabel pdiffusion 863 583 864 584 0 Cellno = 432
rlabel pdiffusion 723 643 724 644 0 Cellno = 433
rlabel pdiffusion 383 303 384 304 0 Cellno = 434
rlabel pdiffusion 423 723 424 724 0 Cellno = 435
rlabel pdiffusion 303 683 304 684 0 Cellno = 436
rlabel pdiffusion 623 663 624 664 0 Cellno = 437
rlabel pdiffusion 703 523 704 524 0 Cellno = 438
rlabel pdiffusion 323 763 324 764 0 Cellno = 439
rlabel pdiffusion 483 783 484 784 0 Cellno = 440
rlabel pdiffusion 703 643 704 644 0 Cellno = 441
rlabel pdiffusion 583 523 584 524 0 Cellno = 442
rlabel pdiffusion 603 523 604 524 0 Cellno = 443
rlabel pdiffusion 463 483 464 484 0 Cellno = 444
rlabel pdiffusion 603 683 604 684 0 Cellno = 445
rlabel pdiffusion 483 703 484 704 0 Cellno = 446
rlabel pdiffusion 763 643 764 644 0 Cellno = 447
rlabel pdiffusion 423 743 424 744 0 Cellno = 448
rlabel pdiffusion 703 263 704 264 0 Cellno = 449
rlabel pdiffusion 443 743 444 744 0 Cellno = 450
rlabel pdiffusion 383 363 384 364 0 Cellno = 451
rlabel pdiffusion 343 603 344 604 0 Cellno = 452
rlabel pdiffusion 563 623 564 624 0 Cellno = 453
rlabel pdiffusion 643 443 644 444 0 Cellno = 454
rlabel pdiffusion 323 283 324 284 0 Cellno = 455
rlabel pdiffusion 663 363 664 364 0 Cellno = 456
rlabel pdiffusion 303 543 304 544 0 Cellno = 457
rlabel pdiffusion 403 703 404 704 0 Cellno = 458
rlabel pdiffusion 623 483 624 484 0 Cellno = 459
rlabel pdiffusion 543 223 544 224 0 Cellno = 460
rlabel pdiffusion 583 343 584 344 0 Cellno = 461
rlabel pdiffusion 503 703 504 704 0 Cellno = 462
rlabel pdiffusion 483 443 484 444 0 Cellno = 463
rlabel pdiffusion 723 543 724 544 0 Cellno = 464
rlabel pdiffusion 303 623 304 624 0 Cellno = 465
rlabel pdiffusion 863 603 864 604 0 Cellno = 466
rlabel pdiffusion 523 683 524 684 0 Cellno = 467
rlabel pdiffusion 763 543 764 544 0 Cellno = 468
rlabel pdiffusion 223 643 224 644 0 Cellno = 469
rlabel pdiffusion 303 503 304 504 0 Cellno = 470
rlabel pdiffusion 403 283 404 284 0 Cellno = 471
rlabel pdiffusion 443 663 444 664 0 Cellno = 472
rlabel pdiffusion 543 603 544 604 0 Cellno = 473
rlabel pdiffusion 363 543 364 544 0 Cellno = 474
rlabel pdiffusion 343 803 344 804 0 Cellno = 475
rlabel pdiffusion 583 643 584 644 0 Cellno = 476
rlabel pdiffusion 503 343 504 344 0 Cellno = 477
rlabel pdiffusion 203 643 204 644 0 Cellno = 478
rlabel pdiffusion 663 803 664 804 0 Cellno = 479
rlabel pdiffusion 163 483 164 484 0 Cellno = 480
rlabel pdiffusion 303 363 304 364 0 Cellno = 481
rlabel pdiffusion 423 543 424 544 0 Cellno = 482
rlabel pdiffusion 623 543 624 544 0 Cellno = 483
rlabel pdiffusion 463 323 464 324 0 Cellno = 484
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 485
rlabel pdiffusion 523 303 524 304 0 Cellno = 486
rlabel pdiffusion 643 363 644 364 0 Cellno = 487
rlabel pdiffusion 223 543 224 544 0 Cellno = 488
rlabel pdiffusion 403 463 404 464 0 Cellno = 489
rlabel pdiffusion 643 603 644 604 0 Cellno = 490
rlabel pdiffusion 883 563 884 564 0 Cellno = 491
rlabel pdiffusion 343 343 344 344 0 Cellno = 492
rlabel pdiffusion 703 443 704 444 0 Cellno = 493
rlabel pdiffusion 423 783 424 784 0 Cellno = 494
rlabel pdiffusion 363 303 364 304 0 Cellno = 495
rlabel pdiffusion 543 623 544 624 0 Cellno = 496
rlabel pdiffusion 363 403 364 404 0 Cellno = 497
rlabel pdiffusion 263 623 264 624 0 Cellno = 498
rlabel pdiffusion 643 483 644 484 0 Cellno = 499
rlabel pdiffusion 643 643 644 644 0 Cellno = 500
rlabel pdiffusion 403 503 404 504 0 Cellno = 501
rlabel pdiffusion 583 743 584 744 0 Cellno = 502
rlabel pdiffusion 143 483 144 484 0 Cellno = 503
rlabel pdiffusion 663 743 664 744 0 Cellno = 504
rlabel pdiffusion 403 843 404 844 0 Cellno = 505
rlabel pdiffusion 383 223 384 224 0 Cellno = 506
rlabel pdiffusion 343 643 344 644 0 Cellno = 507
rlabel pdiffusion 203 423 204 424 0 Cellno = 508
rlabel pdiffusion 763 563 764 564 0 Cellno = 509
rlabel pdiffusion 303 283 304 284 0 Cellno = 510
rlabel pdiffusion 183 623 184 624 0 Cellno = 511
rlabel pdiffusion 423 523 424 524 0 Cellno = 512
rlabel pdiffusion 543 343 544 344 0 Cellno = 513
rlabel pdiffusion 643 383 644 384 0 Cellno = 514
rlabel pdiffusion 803 583 804 584 0 Cellno = 515
rlabel pdiffusion 243 603 244 604 0 Cellno = 516
rlabel pdiffusion 123 563 124 564 0 Cellno = 517
rlabel pdiffusion 803 483 804 484 0 Cellno = 518
rlabel pdiffusion 623 583 624 584 0 Cellno = 519
rlabel pdiffusion 783 563 784 564 0 Cellno = 520
rlabel pdiffusion 843 483 844 484 0 Cellno = 521
rlabel pdiffusion 603 483 604 484 0 Cellno = 522
rlabel pdiffusion 523 803 524 804 0 Cellno = 523
rlabel pdiffusion 483 203 484 204 0 Cellno = 524
rlabel pdiffusion 563 203 564 204 0 Cellno = 525
rlabel pdiffusion 723 403 724 404 0 Cellno = 526
rlabel pdiffusion 283 423 284 424 0 Cellno = 527
rlabel pdiffusion 823 423 824 424 0 Cellno = 528
rlabel pdiffusion 603 243 604 244 0 Cellno = 529
rlabel pdiffusion 623 343 624 344 0 Cellno = 530
rlabel pdiffusion 583 183 584 184 0 Cellno = 531
rlabel pdiffusion 723 623 724 624 0 Cellno = 532
rlabel pdiffusion 463 363 464 364 0 Cellno = 533
rlabel pdiffusion 463 383 464 384 0 Cellno = 534
rlabel pdiffusion 783 403 784 404 0 Cellno = 535
rlabel pdiffusion 603 583 604 584 0 Cellno = 536
rlabel pdiffusion 763 343 764 344 0 Cellno = 537
rlabel pdiffusion 623 603 624 604 0 Cellno = 538
rlabel pdiffusion 563 823 564 824 0 Cellno = 539
rlabel pdiffusion 483 683 484 684 0 Cellno = 540
rlabel pdiffusion 343 523 344 524 0 Cellno = 541
rlabel pdiffusion 183 443 184 444 0 Cellno = 542
rlabel pdiffusion 783 583 784 584 0 Cellno = 543
rlabel pdiffusion 643 683 644 684 0 Cellno = 544
rlabel pdiffusion 703 323 704 324 0 Cellno = 545
rlabel pdiffusion 343 423 344 424 0 Cellno = 546
rlabel pdiffusion 843 603 844 604 0 Cellno = 547
rlabel pdiffusion 303 643 304 644 0 Cellno = 548
rlabel pdiffusion 503 643 504 644 0 Cellno = 549
rlabel pdiffusion 443 523 444 524 0 Cellno = 550
rlabel pdiffusion 323 563 324 564 0 Cellno = 551
rlabel pdiffusion 483 383 484 384 0 Cellno = 552
rlabel pdiffusion 703 483 704 484 0 Cellno = 553
rlabel pdiffusion 383 443 384 444 0 Cellno = 554
rlabel pdiffusion 463 243 464 244 0 Cellno = 555
rlabel pdiffusion 403 363 404 364 0 Cellno = 556
rlabel pdiffusion 603 723 604 724 0 Cellno = 557
rlabel pdiffusion 463 703 464 704 0 Cellno = 558
rlabel pdiffusion 483 563 484 564 0 Cellno = 559
rlabel pdiffusion 663 763 664 764 0 Cellno = 560
rlabel pdiffusion 383 743 384 744 0 Cellno = 561
rlabel pdiffusion 683 763 684 764 0 Cellno = 562
rlabel pdiffusion 643 243 644 244 0 Cellno = 563
rlabel pdiffusion 743 503 744 504 0 Cellno = 564
rlabel pdiffusion 383 703 384 704 0 Cellno = 565
rlabel pdiffusion 383 583 384 584 0 Cellno = 566
rlabel pdiffusion 723 343 724 344 0 Cellno = 567
rlabel pdiffusion 403 183 404 184 0 Cellno = 568
rlabel pdiffusion 383 563 384 564 0 Cellno = 569
rlabel pdiffusion 523 323 524 324 0 Cellno = 570
rlabel pdiffusion 683 303 684 304 0 Cellno = 571
rlabel pdiffusion 663 263 664 264 0 Cellno = 572
rlabel pdiffusion 463 203 464 204 0 Cellno = 573
rlabel pdiffusion 223 623 224 624 0 Cellno = 574
rlabel pdiffusion 383 823 384 824 0 Cellno = 575
rlabel pdiffusion 623 643 624 644 0 Cellno = 576
rlabel pdiffusion 423 443 424 444 0 Cellno = 577
rlabel pdiffusion 323 523 324 524 0 Cellno = 578
rlabel pdiffusion 403 583 404 584 0 Cellno = 579
rlabel pdiffusion 383 803 384 804 0 Cellno = 580
rlabel pdiffusion 603 603 604 604 0 Cellno = 581
rlabel pdiffusion 543 743 544 744 0 Cellno = 582
rlabel pdiffusion 483 623 484 624 0 Cellno = 583
rlabel pdiffusion 803 523 804 524 0 Cellno = 584
rlabel pdiffusion 563 683 564 684 0 Cellno = 585
rlabel pdiffusion 583 623 584 624 0 Cellno = 586
rlabel pdiffusion 243 403 244 404 0 Cellno = 587
rlabel pdiffusion 603 363 604 364 0 Cellno = 588
rlabel pdiffusion 523 883 524 884 0 Cellno = 589
rlabel pdiffusion 543 383 544 384 0 Cellno = 590
rlabel pdiffusion 223 583 224 584 0 Cellno = 591
rlabel pdiffusion 683 743 684 744 0 Cellno = 592
rlabel pdiffusion 403 483 404 484 0 Cellno = 593
rlabel pdiffusion 763 623 764 624 0 Cellno = 594
rlabel pdiffusion 603 763 604 764 0 Cellno = 595
rlabel pdiffusion 603 663 604 664 0 Cellno = 596
rlabel pdiffusion 463 763 464 764 0 Cellno = 597
rlabel pdiffusion 603 323 604 324 0 Cellno = 598
rlabel pdiffusion 703 383 704 384 0 Cellno = 599
rlabel pdiffusion 703 723 704 724 0 Cellno = 600
rlabel pdiffusion 683 783 684 784 0 Cellno = 601
rlabel pdiffusion 543 723 544 724 0 Cellno = 602
rlabel pdiffusion 283 663 284 664 0 Cellno = 603
rlabel pdiffusion 763 443 764 444 0 Cellno = 604
rlabel pdiffusion 503 503 504 504 0 Cellno = 605
rlabel pdiffusion 243 463 244 464 0 Cellno = 606
rlabel pdiffusion 323 403 324 404 0 Cellno = 607
rlabel pdiffusion 543 863 544 864 0 Cellno = 608
rlabel pdiffusion 263 423 264 424 0 Cellno = 609
rlabel pdiffusion 683 623 684 624 0 Cellno = 610
rlabel pdiffusion 323 303 324 304 0 Cellno = 611
rlabel pdiffusion 643 663 644 664 0 Cellno = 612
rlabel pdiffusion 663 723 664 724 0 Cellno = 613
rlabel pdiffusion 583 503 584 504 0 Cellno = 614
rlabel pdiffusion 443 483 444 484 0 Cellno = 615
rlabel pdiffusion 683 803 684 804 0 Cellno = 616
rlabel pdiffusion 623 363 624 364 0 Cellno = 617
rlabel pdiffusion 503 483 504 484 0 Cellno = 618
rlabel pdiffusion 283 703 284 704 0 Cellno = 619
rlabel pdiffusion 203 603 204 604 0 Cellno = 620
rlabel pdiffusion 763 683 764 684 0 Cellno = 621
rlabel pdiffusion 583 543 584 544 0 Cellno = 622
rlabel pdiffusion 123 543 124 544 0 Cellno = 623
rlabel pdiffusion 183 603 184 604 0 Cellno = 624
rlabel pdiffusion 523 383 524 384 0 Cellno = 625
rlabel pdiffusion 503 443 504 444 0 Cellno = 626
rlabel pdiffusion 343 283 344 284 0 Cellno = 627
rlabel pdiffusion 443 423 444 424 0 Cellno = 628
rlabel pdiffusion 743 543 744 544 0 Cellno = 629
rlabel pdiffusion 543 883 544 884 0 Cellno = 630
rlabel pdiffusion 463 283 464 284 0 Cellno = 631
rlabel pdiffusion 383 543 384 544 0 Cellno = 632
rlabel pdiffusion 683 543 684 544 0 Cellno = 633
rlabel pdiffusion 503 303 504 304 0 Cellno = 634
rlabel pdiffusion 363 323 364 324 0 Cellno = 635
rlabel pdiffusion 523 343 524 344 0 Cellno = 636
rlabel pdiffusion 683 323 684 324 0 Cellno = 637
rlabel pdiffusion 543 703 544 704 0 Cellno = 638
rlabel pdiffusion 423 623 424 624 0 Cellno = 639
rlabel pdiffusion 663 563 664 564 0 Cellno = 640
rlabel pdiffusion 543 303 544 304 0 Cellno = 641
rlabel pdiffusion 543 803 544 804 0 Cellno = 642
rlabel pdiffusion 303 463 304 464 0 Cellno = 643
rlabel pdiffusion 583 603 584 604 0 Cellno = 644
rlabel pdiffusion 383 783 384 784 0 Cellno = 645
rlabel pdiffusion 483 483 484 484 0 Cellno = 646
rlabel pdiffusion 403 403 404 404 0 Cellno = 647
rlabel pdiffusion 583 303 584 304 0 Cellno = 648
rlabel pdiffusion 663 423 664 424 0 Cellno = 649
rlabel pdiffusion 203 403 204 404 0 Cellno = 650
rlabel pdiffusion 523 243 524 244 0 Cellno = 651
rlabel pdiffusion 343 663 344 664 0 Cellno = 652
rlabel pdiffusion 803 663 804 664 0 Cellno = 653
rlabel pdiffusion 303 523 304 524 0 Cellno = 654
rlabel pdiffusion 663 303 664 304 0 Cellno = 655
rlabel pdiffusion 603 503 604 504 0 Cellno = 656
rlabel pdiffusion 343 243 344 244 0 Cellno = 657
rlabel pdiffusion 743 423 744 424 0 Cellno = 658
rlabel pdiffusion 583 863 584 864 0 Cellno = 659
rlabel pdiffusion 203 463 204 464 0 Cellno = 660
rlabel pdiffusion 723 383 724 384 0 Cellno = 661
rlabel pdiffusion 423 763 424 764 0 Cellno = 662
rlabel pdiffusion 643 763 644 764 0 Cellno = 663
rlabel pdiffusion 583 383 584 384 0 Cellno = 664
rlabel pdiffusion 563 843 564 844 0 Cellno = 665
rlabel pdiffusion 383 623 384 624 0 Cellno = 666
rlabel pdiffusion 683 463 684 464 0 Cellno = 667
rlabel pdiffusion 463 563 464 564 0 Cellno = 668
rlabel pdiffusion 623 323 624 324 0 Cellno = 669
rlabel pdiffusion 503 363 504 364 0 Cellno = 670
rlabel pdiffusion 603 303 604 304 0 Cellno = 671
rlabel pdiffusion 443 403 444 404 0 Cellno = 672
rlabel pdiffusion 403 723 404 724 0 Cellno = 673
rlabel pdiffusion 883 583 884 584 0 Cellno = 674
rlabel pdiffusion 323 743 324 744 0 Cellno = 675
rlabel pdiffusion 583 843 584 844 0 Cellno = 676
rlabel pdiffusion 523 483 524 484 0 Cellno = 677
rlabel pdiffusion 303 763 304 764 0 Cellno = 678
rlabel pdiffusion 843 523 844 524 0 Cellno = 679
rlabel pdiffusion 403 203 404 204 0 Cellno = 680
rlabel pdiffusion 563 383 564 384 0 Cellno = 681
rlabel pdiffusion 363 243 364 244 0 Cellno = 682
rlabel pdiffusion 383 503 384 504 0 Cellno = 683
rlabel pdiffusion 563 523 564 524 0 Cellno = 684
rlabel pdiffusion 163 643 164 644 0 Cellno = 685
rlabel pdiffusion 583 463 584 464 0 Cellno = 686
rlabel pdiffusion 483 503 484 504 0 Cellno = 687
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 688
rlabel pdiffusion 663 683 664 684 0 Cellno = 689
rlabel pdiffusion 483 603 484 604 0 Cellno = 690
rlabel pdiffusion 243 723 244 724 0 Cellno = 691
rlabel pdiffusion 343 363 344 364 0 Cellno = 692
rlabel pdiffusion 363 643 364 644 0 Cellno = 693
rlabel pdiffusion 403 683 404 684 0 Cellno = 694
rlabel pdiffusion 583 363 584 364 0 Cellno = 695
rlabel pdiffusion 623 283 624 284 0 Cellno = 696
rlabel pdiffusion 603 183 604 184 0 Cellno = 697
rlabel pdiffusion 683 643 684 644 0 Cellno = 698
rlabel pdiffusion 503 163 504 164 0 Cellno = 699
rlabel pdiffusion 563 343 564 344 0 Cellno = 700
rlabel pdiffusion 683 343 684 344 0 Cellno = 701
rlabel pdiffusion 523 903 524 904 0 Cellno = 702
rlabel pdiffusion 583 283 584 284 0 Cellno = 703
rlabel pdiffusion 563 783 564 784 0 Cellno = 704
rlabel pdiffusion 403 383 404 384 0 Cellno = 705
rlabel pdiffusion 283 363 284 364 0 Cellno = 706
rlabel pdiffusion 443 643 444 644 0 Cellno = 707
rlabel pdiffusion 563 183 564 184 0 Cellno = 708
rlabel pdiffusion 783 463 784 464 0 Cellno = 709
rlabel pdiffusion 863 443 864 444 0 Cellno = 710
rlabel pdiffusion 783 603 784 604 0 Cellno = 711
rlabel pdiffusion 363 463 364 464 0 Cellno = 712
rlabel pdiffusion 403 523 404 524 0 Cellno = 713
rlabel pdiffusion 743 343 744 344 0 Cellno = 714
rlabel pdiffusion 823 543 824 544 0 Cellno = 715
rlabel pdiffusion 443 263 444 264 0 Cellno = 716
rlabel pdiffusion 343 463 344 464 0 Cellno = 717
rlabel pdiffusion 663 403 664 404 0 Cellno = 718
rlabel pdiffusion 563 563 564 564 0 Cellno = 719
rlabel pdiffusion 603 263 604 264 0 Cellno = 720
rlabel pdiffusion 783 483 784 484 0 Cellno = 721
rlabel pdiffusion 443 223 444 224 0 Cellno = 722
rlabel pdiffusion 203 563 204 564 0 Cellno = 723
rlabel pdiffusion 183 463 184 464 0 Cellno = 724
rlabel pdiffusion 303 783 304 784 0 Cellno = 725
rlabel pdiffusion 663 703 664 704 0 Cellno = 726
rlabel pdiffusion 603 383 604 384 0 Cellno = 727
rlabel pdiffusion 623 243 624 244 0 Cellno = 728
rlabel pdiffusion 723 703 724 704 0 Cellno = 729
rlabel pdiffusion 423 303 424 304 0 Cellno = 730
rlabel pdiffusion 183 403 184 404 0 Cellno = 731
rlabel pdiffusion 423 243 424 244 0 Cellno = 732
rlabel pdiffusion 523 503 524 504 0 Cellno = 733
rlabel pdiffusion 683 423 684 424 0 Cellno = 734
rlabel pdiffusion 363 483 364 484 0 Cellno = 735
rlabel pdiffusion 763 583 764 584 0 Cellno = 736
rlabel pdiffusion 603 643 604 644 0 Cellno = 737
rlabel pdiffusion 303 403 304 404 0 Cellno = 738
rlabel pdiffusion 203 483 204 484 0 Cellno = 739
rlabel pdiffusion 663 483 664 484 0 Cellno = 740
rlabel pdiffusion 743 563 744 564 0 Cellno = 741
rlabel pdiffusion 723 603 724 604 0 Cellno = 742
rlabel pdiffusion 643 743 644 744 0 Cellno = 743
rlabel pdiffusion 303 343 304 344 0 Cellno = 744
rlabel pdiffusion 723 323 724 324 0 Cellno = 745
rlabel pdiffusion 243 743 244 744 0 Cellno = 746
rlabel pdiffusion 483 883 484 884 0 Cellno = 747
rlabel pdiffusion 563 443 564 444 0 Cellno = 748
rlabel pdiffusion 483 363 484 364 0 Cellno = 749
rlabel pdiffusion 603 543 604 544 0 Cellno = 750
rlabel pdiffusion 663 523 664 524 0 Cellno = 751
rlabel pdiffusion 363 363 364 364 0 Cellno = 752
rlabel pdiffusion 223 383 224 384 0 Cellno = 753
rlabel pdiffusion 823 623 824 624 0 Cellno = 754
rlabel pdiffusion 683 283 684 284 0 Cellno = 755
rlabel pdiffusion 363 683 364 684 0 Cellno = 756
rlabel pdiffusion 363 663 364 664 0 Cellno = 757
rlabel pdiffusion 163 463 164 464 0 Cellno = 758
rlabel pdiffusion 483 523 484 524 0 Cellno = 759
rlabel pdiffusion 363 503 364 504 0 Cellno = 760
rlabel pdiffusion 543 783 544 784 0 Cellno = 761
rlabel pdiffusion 563 123 564 124 0 Cellno = 762
rlabel pdiffusion 743 623 744 624 0 Cellno = 763
rlabel pdiffusion 543 363 544 364 0 Cellno = 764
rlabel pdiffusion 323 443 324 444 0 Cellno = 765
rlabel pdiffusion 663 463 664 464 0 Cellno = 766
rlabel pdiffusion 583 243 584 244 0 Cellno = 767
rlabel pdiffusion 463 823 464 824 0 Cellno = 768
rlabel pdiffusion 623 743 624 744 0 Cellno = 769
rlabel pdiffusion 663 663 664 664 0 Cellno = 770
rlabel pdiffusion 503 323 504 324 0 Cellno = 771
rlabel pdiffusion 703 463 704 464 0 Cellno = 772
rlabel pdiffusion 663 603 664 604 0 Cellno = 773
rlabel pdiffusion 443 703 444 704 0 Cellno = 774
rlabel pdiffusion 243 323 244 324 0 Cellno = 775
rlabel pdiffusion 323 663 324 664 0 Cellno = 776
rlabel pdiffusion 363 723 364 724 0 Cellno = 777
rlabel pdiffusion 403 663 404 664 0 Cellno = 778
rlabel pdiffusion 643 823 644 824 0 Cellno = 779
rlabel pdiffusion 243 703 244 704 0 Cellno = 780
rlabel pdiffusion 623 803 624 804 0 Cellno = 781
rlabel pdiffusion 263 483 264 484 0 Cellno = 782
rlabel pdiffusion 743 463 744 464 0 Cellno = 783
rlabel pdiffusion 683 703 684 704 0 Cellno = 784
rlabel pdiffusion 523 723 524 724 0 Cellno = 785
rlabel pdiffusion 603 343 604 344 0 Cellno = 786
rlabel pdiffusion 443 863 444 864 0 Cellno = 787
rlabel pdiffusion 563 483 564 484 0 Cellno = 788
rlabel pdiffusion 683 263 684 264 0 Cellno = 789
rlabel pdiffusion 483 403 484 404 0 Cellno = 790
rlabel pdiffusion 723 463 724 464 0 Cellno = 791
rlabel pdiffusion 383 243 384 244 0 Cellno = 792
rlabel pdiffusion 443 683 444 684 0 Cellno = 793
rlabel pdiffusion 403 743 404 744 0 Cellno = 794
rlabel pdiffusion 643 423 644 424 0 Cellno = 795
rlabel pdiffusion 283 523 284 524 0 Cellno = 796
rlabel pdiffusion 703 563 704 564 0 Cellno = 797
rlabel pdiffusion 343 623 344 624 0 Cellno = 798
rlabel pdiffusion 523 443 524 444 0 Cellno = 799
rlabel pdiffusion 543 163 544 164 0 Cellno = 800
rlabel pdiffusion 443 343 444 344 0 Cellno = 801
rlabel pdiffusion 803 563 804 564 0 Cellno = 802
rlabel pdiffusion 483 823 484 824 0 Cellno = 803
rlabel pdiffusion 243 623 244 624 0 Cellno = 804
rlabel pdiffusion 323 783 324 784 0 Cellno = 805
rlabel pdiffusion 363 623 364 624 0 Cellno = 806
rlabel pdiffusion 703 763 704 764 0 Cellno = 807
rlabel pdiffusion 423 583 424 584 0 Cellno = 808
rlabel pdiffusion 683 663 684 664 0 Cellno = 809
rlabel pdiffusion 323 263 324 264 0 Cellno = 810
rlabel pdiffusion 803 423 804 424 0 Cellno = 811
rlabel pdiffusion 323 463 324 464 0 Cellno = 812
rlabel pdiffusion 703 363 704 364 0 Cellno = 813
rlabel pdiffusion 603 563 604 564 0 Cellno = 814
rlabel pdiffusion 243 583 244 584 0 Cellno = 815
rlabel pdiffusion 743 643 744 644 0 Cellno = 816
rlabel pdiffusion 743 403 744 404 0 Cellno = 817
rlabel pdiffusion 663 223 664 224 0 Cellno = 818
rlabel pdiffusion 103 523 104 524 0 Cellno = 819
rlabel pdiffusion 363 523 364 524 0 Cellno = 820
rlabel pdiffusion 423 323 424 324 0 Cellno = 821
rlabel pdiffusion 503 723 504 724 0 Cellno = 822
rlabel pdiffusion 743 383 744 384 0 Cellno = 823
rlabel pdiffusion 223 683 224 684 0 Cellno = 824
rlabel pdiffusion 423 363 424 364 0 Cellno = 825
rlabel pdiffusion 263 523 264 524 0 Cellno = 826
rlabel pdiffusion 783 423 784 424 0 Cellno = 827
rlabel pdiffusion 383 643 384 644 0 Cellno = 828
rlabel pdiffusion 523 543 524 544 0 Cellno = 829
rlabel pdiffusion 723 583 724 584 0 Cellno = 830
rlabel pdiffusion 443 463 444 464 0 Cellno = 831
rlabel pdiffusion 663 383 664 384 0 Cellno = 832
rlabel pdiffusion 423 263 424 264 0 Cellno = 833
rlabel pdiffusion 523 703 524 704 0 Cellno = 834
rlabel pdiffusion 683 483 684 484 0 Cellno = 835
rlabel pdiffusion 683 443 684 444 0 Cellno = 836
rlabel pdiffusion 363 563 364 564 0 Cellno = 837
rlabel pdiffusion 603 223 604 224 0 Cellno = 838
rlabel pdiffusion 523 783 524 784 0 Cellno = 839
rlabel pdiffusion 263 683 264 684 0 Cellno = 840
rlabel pdiffusion 543 443 544 444 0 Cellno = 841
rlabel pdiffusion 323 703 324 704 0 Cellno = 842
rlabel pdiffusion 763 383 764 384 0 Cellno = 843
rlabel pdiffusion 423 663 424 664 0 Cellno = 844
rlabel pdiffusion 223 443 224 444 0 Cellno = 845
rlabel pdiffusion 363 423 364 424 0 Cellno = 846
rlabel pdiffusion 783 663 784 664 0 Cellno = 847
rlabel pdiffusion 463 803 464 804 0 Cellno = 848
rlabel pdiffusion 723 663 724 664 0 Cellno = 849
rlabel pdiffusion 563 363 564 364 0 Cellno = 850
rlabel pdiffusion 603 283 604 284 0 Cellno = 851
rlabel pdiffusion 383 463 384 464 0 Cellno = 852
rlabel pdiffusion 583 403 584 404 0 Cellno = 853
rlabel pdiffusion 523 263 524 264 0 Cellno = 854
rlabel pdiffusion 623 303 624 304 0 Cellno = 855
rlabel pdiffusion 283 463 284 464 0 Cellno = 856
rlabel pdiffusion 303 443 304 444 0 Cellno = 857
rlabel pdiffusion 503 203 504 204 0 Cellno = 858
rlabel pdiffusion 143 643 144 644 0 Cellno = 859
rlabel pdiffusion 643 623 644 624 0 Cellno = 860
rlabel pdiffusion 403 343 404 344 0 Cellno = 861
rlabel pdiffusion 883 543 884 544 0 Cellno = 862
rlabel pdiffusion 763 523 764 524 0 Cellno = 863
rlabel pdiffusion 423 463 424 464 0 Cellno = 864
rlabel pdiffusion 483 423 484 424 0 Cellno = 865
rlabel pdiffusion 523 843 524 844 0 Cellno = 866
rlabel pdiffusion 543 663 544 664 0 Cellno = 867
rlabel pdiffusion 463 603 464 604 0 Cellno = 868
rlabel pdiffusion 463 503 464 504 0 Cellno = 869
rlabel pdiffusion 783 503 784 504 0 Cellno = 870
rlabel pdiffusion 343 763 344 764 0 Cellno = 871
rlabel pdiffusion 263 403 264 404 0 Cellno = 872
rlabel pdiffusion 443 283 444 284 0 Cellno = 873
rlabel pdiffusion 683 183 684 184 0 Cellno = 874
rlabel pdiffusion 223 503 224 504 0 Cellno = 875
rlabel pdiffusion 623 843 624 844 0 Cellno = 876
rlabel pdiffusion 543 243 544 244 0 Cellno = 877
rlabel pdiffusion 363 383 364 384 0 Cellno = 878
rlabel pdiffusion 723 483 724 484 0 Cellno = 879
rlabel pdiffusion 283 623 284 624 0 Cellno = 880
rlabel pdiffusion 243 343 244 344 0 Cellno = 881
rlabel pdiffusion 363 743 364 744 0 Cellno = 882
rlabel pdiffusion 383 323 384 324 0 Cellno = 883
rlabel pdiffusion 383 383 384 384 0 Cellno = 884
rlabel pdiffusion 203 583 204 584 0 Cellno = 885
rlabel pdiffusion 403 243 404 244 0 Cellno = 886
rlabel pdiffusion 243 563 244 564 0 Cellno = 887
rlabel pdiffusion 723 523 724 524 0 Cellno = 888
rlabel pdiffusion 663 643 664 644 0 Cellno = 889
rlabel pdiffusion 303 603 304 604 0 Cellno = 890
rlabel pdiffusion 503 743 504 744 0 Cellno = 891
rlabel pdiffusion 603 203 604 204 0 Cellno = 892
rlabel pdiffusion 583 883 584 884 0 Cellno = 893
rlabel pdiffusion 183 503 184 504 0 Cellno = 894
rlabel pdiffusion 583 663 584 664 0 Cellno = 895
rlabel pdiffusion 663 443 664 444 0 Cellno = 896
rlabel pdiffusion 523 463 524 464 0 Cellno = 897
rlabel pdiffusion 463 743 464 744 0 Cellno = 898
rlabel pdiffusion 443 203 444 204 0 Cellno = 899
rlabel pdiffusion 863 563 864 564 0 Cellno = 900
rlabel pdiffusion 303 303 304 304 0 Cellno = 901
rlabel pdiffusion 303 663 304 664 0 Cellno = 902
rlabel pdiffusion 763 403 764 404 0 Cellno = 903
rlabel pdiffusion 343 483 344 484 0 Cellno = 904
rlabel pdiffusion 483 183 484 184 0 Cellno = 905
rlabel pdiffusion 243 523 244 524 0 Cellno = 906
rlabel pdiffusion 643 723 644 724 0 Cellno = 907
rlabel pdiffusion 443 323 444 324 0 Cellno = 908
rlabel pdiffusion 803 543 804 544 0 Cellno = 909
rlabel pdiffusion 343 543 344 544 0 Cellno = 910
rlabel pdiffusion 543 283 544 284 0 Cellno = 911
rlabel pdiffusion 703 403 704 404 0 Cellno = 912
rlabel pdiffusion 543 583 544 584 0 Cellno = 913
rlabel pdiffusion 323 803 324 804 0 Cellno = 914
rlabel pdiffusion 343 503 344 504 0 Cellno = 915
rlabel pdiffusion 543 683 544 684 0 Cellno = 916
rlabel pdiffusion 563 703 564 704 0 Cellno = 917
rlabel pdiffusion 723 303 724 304 0 Cellno = 918
rlabel pdiffusion 563 223 564 224 0 Cellno = 919
rlabel pdiffusion 423 223 424 224 0 Cellno = 920
rlabel pdiffusion 523 223 524 224 0 Cellno = 921
rlabel pdiffusion 283 383 284 384 0 Cellno = 922
rlabel pdiffusion 763 423 764 424 0 Cellno = 923
rlabel pdiffusion 503 543 504 544 0 Cellno = 924
rlabel pdiffusion 443 563 444 564 0 Cellno = 925
rlabel pdiffusion 523 623 524 624 0 Cellno = 926
rlabel pdiffusion 123 523 124 524 0 Cellno = 927
rlabel pdiffusion 603 703 604 704 0 Cellno = 928
rlabel pdiffusion 883 483 884 484 0 Cellno = 929
rlabel pdiffusion 643 463 644 464 0 Cellno = 930
rlabel pdiffusion 503 823 504 824 0 Cellno = 931
rlabel pdiffusion 503 463 504 464 0 Cellno = 932
rlabel pdiffusion 303 583 304 584 0 Cellno = 933
rlabel pdiffusion 643 283 644 284 0 Cellno = 934
rlabel pdiffusion 403 323 404 324 0 Cellno = 935
rlabel pdiffusion 283 323 284 324 0 Cellno = 936
rlabel pdiffusion 803 363 804 364 0 Cellno = 937
rlabel pdiffusion 623 683 624 684 0 Cellno = 938
rlabel pdiffusion 523 203 524 204 0 Cellno = 939
rlabel pdiffusion 843 563 844 564 0 Cellno = 940
rlabel pdiffusion 443 583 444 584 0 Cellno = 941
rlabel pdiffusion 503 623 504 624 0 Cellno = 942
rlabel pdiffusion 503 563 504 564 0 Cellno = 943
rlabel pdiffusion 283 563 284 564 0 Cellno = 944
rlabel pdiffusion 483 743 484 744 0 Cellno = 945
rlabel pdiffusion 643 403 644 404 0 Cellno = 946
rlabel pdiffusion 583 263 584 264 0 Cellno = 947
rlabel pdiffusion 223 523 224 524 0 Cellno = 948
rlabel pdiffusion 403 783 404 784 0 Cellno = 949
rlabel pdiffusion 503 243 504 244 0 Cellno = 950
rlabel pdiffusion 723 563 724 564 0 Cellno = 951
rlabel pdiffusion 423 183 424 184 0 Cellno = 952
rlabel pdiffusion 243 503 244 504 0 Cellno = 953
rlabel pdiffusion 583 443 584 444 0 Cellno = 954
rlabel pdiffusion 783 523 784 524 0 Cellno = 955
rlabel pdiffusion 683 683 684 684 0 Cellno = 956
rlabel pdiffusion 263 643 264 644 0 Cellno = 957
rlabel pdiffusion 863 523 864 524 0 Cellno = 958
rlabel pdiffusion 543 423 544 424 0 Cellno = 959
rlabel pdiffusion 523 163 524 164 0 Cellno = 960
rlabel pdiffusion 563 883 564 884 0 Cellno = 961
rlabel pdiffusion 323 423 324 424 0 Cellno = 962
rlabel pdiffusion 543 523 544 524 0 Cellno = 963
rlabel pdiffusion 583 723 584 724 0 Cellno = 964
rlabel pdiffusion 203 683 204 684 0 Cellno = 965
rlabel pdiffusion 363 583 364 584 0 Cellno = 966
rlabel pdiffusion 623 403 624 404 0 Cellno = 967
rlabel pdiffusion 563 403 564 404 0 Cellno = 968
rlabel pdiffusion 563 263 564 264 0 Cellno = 969
rlabel pdiffusion 763 603 764 604 0 Cellno = 970
rlabel pdiffusion 483 263 484 264 0 Cellno = 971
rlabel pdiffusion 623 763 624 764 0 Cellno = 972
rlabel pdiffusion 763 463 764 464 0 Cellno = 973
rlabel pdiffusion 623 563 624 564 0 Cellno = 974
rlabel pdiffusion 783 703 784 704 0 Cellno = 975
rlabel pdiffusion 583 583 584 584 0 Cellno = 976
rlabel pdiffusion 463 583 464 584 0 Cellno = 977
rlabel pdiffusion 583 423 584 424 0 Cellno = 978
rlabel pdiffusion 663 783 664 784 0 Cellno = 979
rlabel pdiffusion 823 443 824 444 0 Cellno = 980
rlabel pdiffusion 503 283 504 284 0 Cellno = 981
rlabel pdiffusion 563 463 564 464 0 Cellno = 982
rlabel pdiffusion 163 403 164 404 0 Cellno = 983
rlabel pdiffusion 583 563 584 564 0 Cellno = 984
rlabel pdiffusion 583 703 584 704 0 Cellno = 985
rlabel pdiffusion 823 503 824 504 0 Cellno = 986
rlabel pdiffusion 723 743 724 744 0 Cellno = 987
rlabel pdiffusion 443 763 444 764 0 Cellno = 988
rlabel pdiffusion 763 323 764 324 0 Cellno = 989
rlabel pdiffusion 343 703 344 704 0 Cellno = 990
rlabel pdiffusion 723 363 724 364 0 Cellno = 991
rlabel pdiffusion 703 703 704 704 0 Cellno = 992
rlabel pdiffusion 523 763 524 764 0 Cellno = 993
rlabel pdiffusion 523 363 524 364 0 Cellno = 994
rlabel pdiffusion 423 563 424 564 0 Cellno = 995
rlabel pdiffusion 163 543 164 544 0 Cellno = 996
rlabel pdiffusion 343 683 344 684 0 Cellno = 997
rlabel pdiffusion 683 363 684 364 0 Cellno = 998
rlabel pdiffusion 223 663 224 664 0 Cellno = 999
rlabel pdiffusion 143 503 144 504 0 Cellno = 1000
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1001
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1002
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1003
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1004
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1005
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1006
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1007
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1008
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1009
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1010
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1011
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1012
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1013
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1014
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1015
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1016
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1017
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1018
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1019
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1020
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1021
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1022
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1023
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1024
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1025
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1026
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1027
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1028
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1029
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1030
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1031
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1032
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1033
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1034
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1035
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1036
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1037
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1038
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1039
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1040
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1041
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1042
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1043
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1044
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1045
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1046
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1047
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1048
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1049
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1050
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1051
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1052
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1053
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1054
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1055
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1056
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1057
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1058
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1059
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1060
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1061
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1062
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1063
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1064
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1065
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1066
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1067
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1068
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1069
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1070
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1071
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1072
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1073
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1074
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1075
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1076
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1077
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1078
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1079
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1080
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1081
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1082
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1083
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1084
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1085
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1086
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1087
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1088
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1089
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1090
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1091
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1092
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1093
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1094
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1095
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1096
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1097
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1098
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1099
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1100
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1101
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1102
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1103
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1104
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1105
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1106
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1107
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1108
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1109
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1110
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1111
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1112
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1113
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1114
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1115
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1116
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1117
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1118
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1119
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1120
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1121
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1122
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1123
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1124
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1125
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1126
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1127
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1128
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1129
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1130
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1131
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1132
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1133
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1134
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1135
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1136
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1137
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1138
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1139
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1140
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1141
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1142
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1143
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1144
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1145
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1146
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1147
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1148
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1149
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1150
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1151
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1152
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1153
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1154
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1155
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1156
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1157
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1158
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1159
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1160
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1161
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1162
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1163
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1164
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1165
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1166
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1167
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1168
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1169
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1170
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1171
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1172
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1173
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1174
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1175
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1176
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1177
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1178
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1179
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1180
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1181
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1182
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1183
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1184
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1185
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1186
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1187
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1188
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1189
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1190
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1191
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1192
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1193
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1194
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1195
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1196
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1197
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1198
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1199
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1200
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1201
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1202
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1203
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1204
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1205
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1206
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1207
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1208
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1209
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1210
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1211
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1212
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1213
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1214
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1215
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1216
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1217
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1218
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1219
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1220
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1221
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1222
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1223
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1224
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1225
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1226
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1227
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1228
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1229
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1230
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1231
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1232
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1233
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1234
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1235
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1236
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1237
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1238
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1239
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1240
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1241
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1242
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1243
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1244
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1245
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1246
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1247
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1248
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1249
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1250
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1251
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1252
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1253
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1254
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1255
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1256
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1257
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1258
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1259
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1260
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1261
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1262
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1263
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1264
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1265
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1266
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1267
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1268
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1269
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1270
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1271
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1272
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1273
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1274
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1275
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1276
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1277
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1278
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1279
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1280
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1281
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1282
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1283
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1284
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1285
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1286
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1287
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1288
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1289
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1290
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1291
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1292
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1293
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1294
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1295
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1296
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1297
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1298
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1299
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1300
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1301
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1302
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1303
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1304
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1305
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1306
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1307
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1308
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1309
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1310
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1311
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1312
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1313
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1314
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1315
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1316
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1317
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1318
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1319
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1320
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1321
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1322
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1323
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1324
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1325
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1326
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1327
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1328
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1329
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1330
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1331
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1332
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1333
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1334
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1335
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1336
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1337
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1338
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1339
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1340
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1341
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1342
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1343
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1344
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1345
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1346
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1347
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1348
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1349
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1350
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1351
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1352
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1353
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1354
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1355
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1356
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1357
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1358
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1359
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1360
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1361
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1362
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1363
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1364
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1365
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1366
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1367
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1368
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1369
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1370
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1371
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1372
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1373
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1374
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1375
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1376
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1377
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1378
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1379
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1380
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1381
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1382
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1383
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1384
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1385
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1386
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1387
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1388
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1389
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1390
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1391
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1392
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1393
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1394
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1395
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1396
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1397
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1398
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1399
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1400
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1401
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1402
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1403
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1404
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1405
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1406
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1407
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1408
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1409
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1410
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1411
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1412
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1413
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1414
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1415
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1416
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1417
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1418
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1419
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1420
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1421
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1422
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1423
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1424
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1425
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1426
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1427
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1428
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1429
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1430
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1431
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1432
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1433
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1434
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1435
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1436
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1437
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1438
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1439
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1440
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1441
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1442
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1443
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1444
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1445
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1446
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1447
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1448
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1449
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1450
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1451
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1452
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1453
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1454
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1455
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1456
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1457
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1458
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1459
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1460
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1461
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1462
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1463
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1464
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1465
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1466
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1467
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1468
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1469
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1470
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1471
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1472
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1473
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1474
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1475
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1476
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1477
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1478
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1479
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1480
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1481
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1482
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1483
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1484
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1485
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1486
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1487
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1488
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1489
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1490
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1491
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1492
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1493
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1494
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1495
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1496
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1497
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1498
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1499
rlabel pdiffusion -17 -17 -16 -16 0 Cellno = 1500
<< end >>
